// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Sep 18 2020 18:21:15

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "SPI" view "INTERFACE"

module SPI (
    ch5_B,
    PWM6,
    ch3_A,
    ch0_B,
    PWM1,
    ch4_B,
    RST,
    PWM0,
    MOSI,
    ch7_B,
    PWM3,
    ch2_B,
    SSEL,
    PWM2,
    MISO,
    ch6_B,
    ch2_A,
    PWM5,
    ch7_A,
    ch6_A,
    ch3_B,
    ch1_A,
    ch0_A,
    SCK,
    PWM4,
    CLK,
    ch5_A,
    ch4_A,
    ch1_B,
    PWM7);

    input ch5_B;
    output PWM6;
    input ch3_A;
    input ch0_B;
    output PWM1;
    input ch4_B;
    input RST;
    output PWM0;
    input MOSI;
    input ch7_B;
    output PWM3;
    input ch2_B;
    input SSEL;
    output PWM2;
    output MISO;
    input ch6_B;
    input ch2_A;
    output PWM5;
    input ch7_A;
    input ch6_A;
    input ch3_B;
    input ch1_A;
    input ch0_A;
    input SCK;
    output PWM4;
    input CLK;
    input ch5_A;
    input ch4_A;
    input ch1_B;
    output PWM7;

    wire N__39370;
    wire N__39369;
    wire N__39368;
    wire N__39361;
    wire N__39360;
    wire N__39359;
    wire N__39352;
    wire N__39351;
    wire N__39350;
    wire N__39343;
    wire N__39342;
    wire N__39341;
    wire N__39334;
    wire N__39333;
    wire N__39332;
    wire N__39325;
    wire N__39324;
    wire N__39323;
    wire N__39316;
    wire N__39315;
    wire N__39314;
    wire N__39307;
    wire N__39306;
    wire N__39305;
    wire N__39298;
    wire N__39297;
    wire N__39296;
    wire N__39289;
    wire N__39288;
    wire N__39287;
    wire N__39280;
    wire N__39279;
    wire N__39278;
    wire N__39271;
    wire N__39270;
    wire N__39269;
    wire N__39262;
    wire N__39261;
    wire N__39260;
    wire N__39253;
    wire N__39252;
    wire N__39251;
    wire N__39244;
    wire N__39243;
    wire N__39242;
    wire N__39235;
    wire N__39234;
    wire N__39233;
    wire N__39226;
    wire N__39225;
    wire N__39224;
    wire N__39217;
    wire N__39216;
    wire N__39215;
    wire N__39208;
    wire N__39207;
    wire N__39206;
    wire N__39199;
    wire N__39198;
    wire N__39197;
    wire N__39190;
    wire N__39189;
    wire N__39188;
    wire N__39181;
    wire N__39180;
    wire N__39179;
    wire N__39172;
    wire N__39171;
    wire N__39170;
    wire N__39163;
    wire N__39162;
    wire N__39161;
    wire N__39154;
    wire N__39153;
    wire N__39152;
    wire N__39145;
    wire N__39144;
    wire N__39143;
    wire N__39136;
    wire N__39135;
    wire N__39134;
    wire N__39127;
    wire N__39126;
    wire N__39125;
    wire N__39118;
    wire N__39117;
    wire N__39116;
    wire N__39109;
    wire N__39108;
    wire N__39107;
    wire N__39090;
    wire N__39087;
    wire N__39084;
    wire N__39081;
    wire N__39078;
    wire N__39075;
    wire N__39072;
    wire N__39069;
    wire N__39066;
    wire N__39065;
    wire N__39064;
    wire N__39057;
    wire N__39056;
    wire N__39055;
    wire N__39054;
    wire N__39053;
    wire N__39050;
    wire N__39049;
    wire N__39048;
    wire N__39047;
    wire N__39046;
    wire N__39037;
    wire N__39036;
    wire N__39035;
    wire N__39034;
    wire N__39031;
    wire N__39024;
    wire N__39021;
    wire N__39018;
    wire N__39011;
    wire N__39006;
    wire N__38997;
    wire N__38994;
    wire N__38993;
    wire N__38988;
    wire N__38985;
    wire N__38984;
    wire N__38983;
    wire N__38982;
    wire N__38979;
    wire N__38972;
    wire N__38967;
    wire N__38966;
    wire N__38965;
    wire N__38962;
    wire N__38957;
    wire N__38952;
    wire N__38951;
    wire N__38948;
    wire N__38947;
    wire N__38946;
    wire N__38943;
    wire N__38938;
    wire N__38937;
    wire N__38934;
    wire N__38933;
    wire N__38932;
    wire N__38929;
    wire N__38926;
    wire N__38923;
    wire N__38920;
    wire N__38917;
    wire N__38914;
    wire N__38913;
    wire N__38912;
    wire N__38911;
    wire N__38910;
    wire N__38905;
    wire N__38902;
    wire N__38901;
    wire N__38900;
    wire N__38893;
    wire N__38890;
    wire N__38887;
    wire N__38884;
    wire N__38883;
    wire N__38880;
    wire N__38879;
    wire N__38878;
    wire N__38877;
    wire N__38872;
    wire N__38869;
    wire N__38866;
    wire N__38865;
    wire N__38864;
    wire N__38857;
    wire N__38852;
    wire N__38847;
    wire N__38842;
    wire N__38837;
    wire N__38834;
    wire N__38831;
    wire N__38828;
    wire N__38825;
    wire N__38818;
    wire N__38805;
    wire N__38802;
    wire N__38799;
    wire N__38798;
    wire N__38797;
    wire N__38796;
    wire N__38795;
    wire N__38794;
    wire N__38793;
    wire N__38790;
    wire N__38787;
    wire N__38782;
    wire N__38777;
    wire N__38774;
    wire N__38763;
    wire N__38762;
    wire N__38761;
    wire N__38760;
    wire N__38759;
    wire N__38758;
    wire N__38755;
    wire N__38752;
    wire N__38747;
    wire N__38744;
    wire N__38741;
    wire N__38738;
    wire N__38735;
    wire N__38724;
    wire N__38723;
    wire N__38722;
    wire N__38721;
    wire N__38720;
    wire N__38719;
    wire N__38718;
    wire N__38717;
    wire N__38716;
    wire N__38715;
    wire N__38714;
    wire N__38713;
    wire N__38712;
    wire N__38711;
    wire N__38710;
    wire N__38709;
    wire N__38708;
    wire N__38707;
    wire N__38706;
    wire N__38705;
    wire N__38704;
    wire N__38703;
    wire N__38702;
    wire N__38701;
    wire N__38700;
    wire N__38699;
    wire N__38698;
    wire N__38697;
    wire N__38696;
    wire N__38695;
    wire N__38694;
    wire N__38693;
    wire N__38692;
    wire N__38691;
    wire N__38690;
    wire N__38689;
    wire N__38688;
    wire N__38687;
    wire N__38686;
    wire N__38685;
    wire N__38684;
    wire N__38683;
    wire N__38682;
    wire N__38681;
    wire N__38680;
    wire N__38679;
    wire N__38678;
    wire N__38677;
    wire N__38676;
    wire N__38675;
    wire N__38674;
    wire N__38673;
    wire N__38672;
    wire N__38671;
    wire N__38670;
    wire N__38669;
    wire N__38668;
    wire N__38667;
    wire N__38666;
    wire N__38665;
    wire N__38664;
    wire N__38663;
    wire N__38662;
    wire N__38661;
    wire N__38660;
    wire N__38659;
    wire N__38658;
    wire N__38657;
    wire N__38656;
    wire N__38655;
    wire N__38654;
    wire N__38653;
    wire N__38652;
    wire N__38651;
    wire N__38650;
    wire N__38649;
    wire N__38648;
    wire N__38647;
    wire N__38646;
    wire N__38645;
    wire N__38644;
    wire N__38643;
    wire N__38642;
    wire N__38641;
    wire N__38640;
    wire N__38639;
    wire N__38638;
    wire N__38637;
    wire N__38636;
    wire N__38635;
    wire N__38634;
    wire N__38633;
    wire N__38632;
    wire N__38631;
    wire N__38630;
    wire N__38629;
    wire N__38628;
    wire N__38627;
    wire N__38626;
    wire N__38625;
    wire N__38624;
    wire N__38623;
    wire N__38622;
    wire N__38621;
    wire N__38620;
    wire N__38619;
    wire N__38618;
    wire N__38617;
    wire N__38616;
    wire N__38615;
    wire N__38614;
    wire N__38613;
    wire N__38612;
    wire N__38611;
    wire N__38610;
    wire N__38609;
    wire N__38608;
    wire N__38607;
    wire N__38606;
    wire N__38605;
    wire N__38604;
    wire N__38603;
    wire N__38602;
    wire N__38601;
    wire N__38600;
    wire N__38599;
    wire N__38598;
    wire N__38597;
    wire N__38596;
    wire N__38595;
    wire N__38594;
    wire N__38593;
    wire N__38592;
    wire N__38591;
    wire N__38590;
    wire N__38589;
    wire N__38588;
    wire N__38587;
    wire N__38586;
    wire N__38585;
    wire N__38584;
    wire N__38583;
    wire N__38582;
    wire N__38581;
    wire N__38580;
    wire N__38579;
    wire N__38578;
    wire N__38577;
    wire N__38576;
    wire N__38575;
    wire N__38574;
    wire N__38573;
    wire N__38572;
    wire N__38571;
    wire N__38570;
    wire N__38569;
    wire N__38568;
    wire N__38567;
    wire N__38566;
    wire N__38565;
    wire N__38564;
    wire N__38563;
    wire N__38562;
    wire N__38561;
    wire N__38560;
    wire N__38559;
    wire N__38558;
    wire N__38557;
    wire N__38556;
    wire N__38555;
    wire N__38554;
    wire N__38553;
    wire N__38552;
    wire N__38551;
    wire N__38550;
    wire N__38549;
    wire N__38548;
    wire N__38547;
    wire N__38546;
    wire N__38545;
    wire N__38544;
    wire N__38543;
    wire N__38542;
    wire N__38541;
    wire N__38172;
    wire N__38169;
    wire N__38166;
    wire N__38163;
    wire N__38160;
    wire N__38159;
    wire N__38158;
    wire N__38157;
    wire N__38156;
    wire N__38155;
    wire N__38154;
    wire N__38153;
    wire N__38152;
    wire N__38149;
    wire N__38146;
    wire N__38143;
    wire N__38140;
    wire N__38139;
    wire N__38138;
    wire N__38137;
    wire N__38132;
    wire N__38129;
    wire N__38126;
    wire N__38123;
    wire N__38118;
    wire N__38115;
    wire N__38114;
    wire N__38113;
    wire N__38110;
    wire N__38107;
    wire N__38104;
    wire N__38101;
    wire N__38100;
    wire N__38097;
    wire N__38096;
    wire N__38095;
    wire N__38094;
    wire N__38091;
    wire N__38088;
    wire N__38085;
    wire N__38080;
    wire N__38077;
    wire N__38074;
    wire N__38067;
    wire N__38064;
    wire N__38061;
    wire N__38058;
    wire N__38055;
    wire N__38052;
    wire N__38049;
    wire N__38042;
    wire N__38037;
    wire N__38030;
    wire N__38013;
    wire N__38010;
    wire N__38007;
    wire N__38004;
    wire N__38001;
    wire N__37998;
    wire N__37995;
    wire N__37992;
    wire N__37989;
    wire N__37986;
    wire N__37985;
    wire N__37984;
    wire N__37977;
    wire N__37974;
    wire N__37971;
    wire N__37968;
    wire N__37965;
    wire N__37962;
    wire N__37961;
    wire N__37960;
    wire N__37957;
    wire N__37954;
    wire N__37951;
    wire N__37946;
    wire N__37941;
    wire N__37938;
    wire N__37935;
    wire N__37932;
    wire N__37929;
    wire N__37926;
    wire N__37923;
    wire N__37920;
    wire N__37917;
    wire N__37914;
    wire N__37911;
    wire N__37908;
    wire N__37905;
    wire N__37902;
    wire N__37899;
    wire N__37896;
    wire N__37895;
    wire N__37890;
    wire N__37887;
    wire N__37886;
    wire N__37885;
    wire N__37884;
    wire N__37881;
    wire N__37878;
    wire N__37873;
    wire N__37868;
    wire N__37863;
    wire N__37860;
    wire N__37857;
    wire N__37854;
    wire N__37851;
    wire N__37848;
    wire N__37845;
    wire N__37842;
    wire N__37839;
    wire N__37836;
    wire N__37833;
    wire N__37830;
    wire N__37827;
    wire N__37824;
    wire N__37821;
    wire N__37818;
    wire N__37815;
    wire N__37812;
    wire N__37811;
    wire N__37810;
    wire N__37807;
    wire N__37802;
    wire N__37799;
    wire N__37794;
    wire N__37791;
    wire N__37788;
    wire N__37787;
    wire N__37784;
    wire N__37783;
    wire N__37780;
    wire N__37777;
    wire N__37774;
    wire N__37767;
    wire N__37764;
    wire N__37763;
    wire N__37762;
    wire N__37761;
    wire N__37760;
    wire N__37759;
    wire N__37756;
    wire N__37749;
    wire N__37748;
    wire N__37745;
    wire N__37744;
    wire N__37743;
    wire N__37742;
    wire N__37741;
    wire N__37738;
    wire N__37737;
    wire N__37734;
    wire N__37731;
    wire N__37728;
    wire N__37725;
    wire N__37722;
    wire N__37719;
    wire N__37716;
    wire N__37713;
    wire N__37712;
    wire N__37709;
    wire N__37708;
    wire N__37705;
    wire N__37704;
    wire N__37703;
    wire N__37702;
    wire N__37701;
    wire N__37694;
    wire N__37689;
    wire N__37686;
    wire N__37681;
    wire N__37678;
    wire N__37675;
    wire N__37672;
    wire N__37669;
    wire N__37666;
    wire N__37663;
    wire N__37660;
    wire N__37657;
    wire N__37654;
    wire N__37647;
    wire N__37640;
    wire N__37637;
    wire N__37634;
    wire N__37617;
    wire N__37614;
    wire N__37613;
    wire N__37612;
    wire N__37609;
    wire N__37606;
    wire N__37603;
    wire N__37600;
    wire N__37595;
    wire N__37592;
    wire N__37589;
    wire N__37586;
    wire N__37583;
    wire N__37578;
    wire N__37575;
    wire N__37572;
    wire N__37569;
    wire N__37566;
    wire N__37565;
    wire N__37564;
    wire N__37563;
    wire N__37562;
    wire N__37561;
    wire N__37560;
    wire N__37559;
    wire N__37558;
    wire N__37557;
    wire N__37556;
    wire N__37553;
    wire N__37550;
    wire N__37547;
    wire N__37544;
    wire N__37541;
    wire N__37538;
    wire N__37537;
    wire N__37534;
    wire N__37531;
    wire N__37528;
    wire N__37525;
    wire N__37522;
    wire N__37521;
    wire N__37514;
    wire N__37513;
    wire N__37512;
    wire N__37511;
    wire N__37508;
    wire N__37507;
    wire N__37506;
    wire N__37505;
    wire N__37504;
    wire N__37503;
    wire N__37502;
    wire N__37499;
    wire N__37496;
    wire N__37493;
    wire N__37486;
    wire N__37483;
    wire N__37480;
    wire N__37477;
    wire N__37474;
    wire N__37469;
    wire N__37466;
    wire N__37463;
    wire N__37456;
    wire N__37449;
    wire N__37444;
    wire N__37439;
    wire N__37434;
    wire N__37427;
    wire N__37410;
    wire N__37407;
    wire N__37404;
    wire N__37401;
    wire N__37398;
    wire N__37395;
    wire N__37394;
    wire N__37389;
    wire N__37388;
    wire N__37387;
    wire N__37386;
    wire N__37385;
    wire N__37382;
    wire N__37381;
    wire N__37380;
    wire N__37379;
    wire N__37378;
    wire N__37375;
    wire N__37374;
    wire N__37371;
    wire N__37366;
    wire N__37363;
    wire N__37360;
    wire N__37357;
    wire N__37352;
    wire N__37351;
    wire N__37348;
    wire N__37345;
    wire N__37344;
    wire N__37341;
    wire N__37338;
    wire N__37333;
    wire N__37332;
    wire N__37327;
    wire N__37324;
    wire N__37323;
    wire N__37322;
    wire N__37317;
    wire N__37314;
    wire N__37313;
    wire N__37312;
    wire N__37307;
    wire N__37304;
    wire N__37301;
    wire N__37296;
    wire N__37293;
    wire N__37290;
    wire N__37285;
    wire N__37280;
    wire N__37263;
    wire N__37260;
    wire N__37257;
    wire N__37254;
    wire N__37251;
    wire N__37250;
    wire N__37247;
    wire N__37246;
    wire N__37245;
    wire N__37244;
    wire N__37243;
    wire N__37242;
    wire N__37241;
    wire N__37240;
    wire N__37237;
    wire N__37234;
    wire N__37231;
    wire N__37228;
    wire N__37225;
    wire N__37224;
    wire N__37221;
    wire N__37218;
    wire N__37215;
    wire N__37212;
    wire N__37211;
    wire N__37210;
    wire N__37207;
    wire N__37202;
    wire N__37197;
    wire N__37194;
    wire N__37191;
    wire N__37186;
    wire N__37183;
    wire N__37180;
    wire N__37177;
    wire N__37174;
    wire N__37171;
    wire N__37168;
    wire N__37165;
    wire N__37160;
    wire N__37155;
    wire N__37152;
    wire N__37137;
    wire N__37136;
    wire N__37135;
    wire N__37134;
    wire N__37133;
    wire N__37132;
    wire N__37131;
    wire N__37130;
    wire N__37129;
    wire N__37128;
    wire N__37125;
    wire N__37122;
    wire N__37119;
    wire N__37116;
    wire N__37115;
    wire N__37112;
    wire N__37109;
    wire N__37106;
    wire N__37103;
    wire N__37100;
    wire N__37099;
    wire N__37096;
    wire N__37093;
    wire N__37090;
    wire N__37087;
    wire N__37084;
    wire N__37081;
    wire N__37078;
    wire N__37075;
    wire N__37072;
    wire N__37067;
    wire N__37064;
    wire N__37061;
    wire N__37060;
    wire N__37055;
    wire N__37050;
    wire N__37047;
    wire N__37038;
    wire N__37033;
    wire N__37030;
    wire N__37017;
    wire N__37014;
    wire N__37013;
    wire N__37012;
    wire N__37009;
    wire N__37006;
    wire N__37003;
    wire N__37000;
    wire N__36995;
    wire N__36992;
    wire N__36989;
    wire N__36984;
    wire N__36981;
    wire N__36980;
    wire N__36977;
    wire N__36974;
    wire N__36973;
    wire N__36970;
    wire N__36967;
    wire N__36964;
    wire N__36961;
    wire N__36958;
    wire N__36955;
    wire N__36948;
    wire N__36945;
    wire N__36942;
    wire N__36939;
    wire N__36936;
    wire N__36933;
    wire N__36932;
    wire N__36929;
    wire N__36926;
    wire N__36925;
    wire N__36920;
    wire N__36917;
    wire N__36916;
    wire N__36913;
    wire N__36910;
    wire N__36907;
    wire N__36906;
    wire N__36899;
    wire N__36896;
    wire N__36893;
    wire N__36890;
    wire N__36887;
    wire N__36884;
    wire N__36881;
    wire N__36878;
    wire N__36873;
    wire N__36872;
    wire N__36871;
    wire N__36868;
    wire N__36865;
    wire N__36862;
    wire N__36859;
    wire N__36856;
    wire N__36853;
    wire N__36850;
    wire N__36847;
    wire N__36844;
    wire N__36841;
    wire N__36838;
    wire N__36831;
    wire N__36828;
    wire N__36827;
    wire N__36824;
    wire N__36821;
    wire N__36818;
    wire N__36817;
    wire N__36814;
    wire N__36811;
    wire N__36808;
    wire N__36805;
    wire N__36800;
    wire N__36795;
    wire N__36792;
    wire N__36789;
    wire N__36786;
    wire N__36783;
    wire N__36780;
    wire N__36777;
    wire N__36776;
    wire N__36773;
    wire N__36770;
    wire N__36767;
    wire N__36766;
    wire N__36763;
    wire N__36760;
    wire N__36757;
    wire N__36750;
    wire N__36747;
    wire N__36746;
    wire N__36743;
    wire N__36740;
    wire N__36739;
    wire N__36736;
    wire N__36733;
    wire N__36730;
    wire N__36727;
    wire N__36722;
    wire N__36719;
    wire N__36716;
    wire N__36711;
    wire N__36708;
    wire N__36705;
    wire N__36702;
    wire N__36699;
    wire N__36696;
    wire N__36693;
    wire N__36690;
    wire N__36687;
    wire N__36684;
    wire N__36681;
    wire N__36678;
    wire N__36675;
    wire N__36672;
    wire N__36669;
    wire N__36666;
    wire N__36663;
    wire N__36660;
    wire N__36657;
    wire N__36654;
    wire N__36651;
    wire N__36648;
    wire N__36645;
    wire N__36642;
    wire N__36639;
    wire N__36636;
    wire N__36633;
    wire N__36630;
    wire N__36629;
    wire N__36626;
    wire N__36623;
    wire N__36618;
    wire N__36617;
    wire N__36616;
    wire N__36613;
    wire N__36610;
    wire N__36607;
    wire N__36604;
    wire N__36597;
    wire N__36596;
    wire N__36595;
    wire N__36592;
    wire N__36589;
    wire N__36586;
    wire N__36581;
    wire N__36576;
    wire N__36575;
    wire N__36574;
    wire N__36569;
    wire N__36566;
    wire N__36563;
    wire N__36558;
    wire N__36557;
    wire N__36556;
    wire N__36553;
    wire N__36550;
    wire N__36547;
    wire N__36544;
    wire N__36537;
    wire N__36534;
    wire N__36531;
    wire N__36528;
    wire N__36525;
    wire N__36522;
    wire N__36521;
    wire N__36518;
    wire N__36515;
    wire N__36514;
    wire N__36513;
    wire N__36512;
    wire N__36507;
    wire N__36504;
    wire N__36503;
    wire N__36502;
    wire N__36501;
    wire N__36498;
    wire N__36495;
    wire N__36494;
    wire N__36489;
    wire N__36488;
    wire N__36487;
    wire N__36486;
    wire N__36485;
    wire N__36484;
    wire N__36483;
    wire N__36480;
    wire N__36477;
    wire N__36474;
    wire N__36471;
    wire N__36468;
    wire N__36465;
    wire N__36462;
    wire N__36451;
    wire N__36448;
    wire N__36445;
    wire N__36442;
    wire N__36439;
    wire N__36438;
    wire N__36435;
    wire N__36430;
    wire N__36427;
    wire N__36424;
    wire N__36421;
    wire N__36418;
    wire N__36415;
    wire N__36412;
    wire N__36409;
    wire N__36402;
    wire N__36397;
    wire N__36384;
    wire N__36381;
    wire N__36378;
    wire N__36377;
    wire N__36376;
    wire N__36373;
    wire N__36372;
    wire N__36371;
    wire N__36370;
    wire N__36369;
    wire N__36368;
    wire N__36367;
    wire N__36366;
    wire N__36363;
    wire N__36362;
    wire N__36359;
    wire N__36348;
    wire N__36347;
    wire N__36346;
    wire N__36345;
    wire N__36342;
    wire N__36339;
    wire N__36336;
    wire N__36333;
    wire N__36332;
    wire N__36329;
    wire N__36326;
    wire N__36323;
    wire N__36320;
    wire N__36317;
    wire N__36314;
    wire N__36311;
    wire N__36308;
    wire N__36305;
    wire N__36302;
    wire N__36299;
    wire N__36296;
    wire N__36293;
    wire N__36290;
    wire N__36285;
    wire N__36284;
    wire N__36281;
    wire N__36278;
    wire N__36271;
    wire N__36266;
    wire N__36263;
    wire N__36260;
    wire N__36257;
    wire N__36254;
    wire N__36251;
    wire N__36246;
    wire N__36239;
    wire N__36236;
    wire N__36225;
    wire N__36222;
    wire N__36219;
    wire N__36218;
    wire N__36217;
    wire N__36212;
    wire N__36209;
    wire N__36206;
    wire N__36201;
    wire N__36200;
    wire N__36197;
    wire N__36196;
    wire N__36193;
    wire N__36190;
    wire N__36187;
    wire N__36184;
    wire N__36181;
    wire N__36174;
    wire N__36171;
    wire N__36168;
    wire N__36167;
    wire N__36166;
    wire N__36165;
    wire N__36164;
    wire N__36161;
    wire N__36160;
    wire N__36159;
    wire N__36158;
    wire N__36157;
    wire N__36154;
    wire N__36151;
    wire N__36150;
    wire N__36149;
    wire N__36146;
    wire N__36143;
    wire N__36142;
    wire N__36139;
    wire N__36136;
    wire N__36135;
    wire N__36134;
    wire N__36133;
    wire N__36130;
    wire N__36127;
    wire N__36124;
    wire N__36121;
    wire N__36118;
    wire N__36115;
    wire N__36112;
    wire N__36109;
    wire N__36106;
    wire N__36103;
    wire N__36098;
    wire N__36095;
    wire N__36090;
    wire N__36089;
    wire N__36084;
    wire N__36081;
    wire N__36076;
    wire N__36073;
    wire N__36070;
    wire N__36065;
    wire N__36062;
    wire N__36055;
    wire N__36052;
    wire N__36049;
    wire N__36046;
    wire N__36037;
    wire N__36030;
    wire N__36021;
    wire N__36018;
    wire N__36015;
    wire N__36014;
    wire N__36013;
    wire N__36012;
    wire N__36011;
    wire N__36010;
    wire N__36007;
    wire N__36006;
    wire N__36005;
    wire N__36004;
    wire N__36003;
    wire N__36002;
    wire N__35999;
    wire N__35998;
    wire N__35995;
    wire N__35994;
    wire N__35993;
    wire N__35990;
    wire N__35987;
    wire N__35978;
    wire N__35975;
    wire N__35974;
    wire N__35973;
    wire N__35970;
    wire N__35967;
    wire N__35964;
    wire N__35961;
    wire N__35958;
    wire N__35955;
    wire N__35952;
    wire N__35949;
    wire N__35944;
    wire N__35941;
    wire N__35938;
    wire N__35935;
    wire N__35930;
    wire N__35927;
    wire N__35924;
    wire N__35919;
    wire N__35916;
    wire N__35911;
    wire N__35906;
    wire N__35903;
    wire N__35900;
    wire N__35897;
    wire N__35892;
    wire N__35887;
    wire N__35882;
    wire N__35871;
    wire N__35868;
    wire N__35865;
    wire N__35862;
    wire N__35861;
    wire N__35858;
    wire N__35855;
    wire N__35854;
    wire N__35853;
    wire N__35848;
    wire N__35845;
    wire N__35842;
    wire N__35839;
    wire N__35832;
    wire N__35831;
    wire N__35830;
    wire N__35829;
    wire N__35828;
    wire N__35827;
    wire N__35826;
    wire N__35825;
    wire N__35824;
    wire N__35821;
    wire N__35818;
    wire N__35815;
    wire N__35812;
    wire N__35809;
    wire N__35806;
    wire N__35803;
    wire N__35800;
    wire N__35797;
    wire N__35796;
    wire N__35795;
    wire N__35794;
    wire N__35793;
    wire N__35790;
    wire N__35789;
    wire N__35788;
    wire N__35787;
    wire N__35786;
    wire N__35785;
    wire N__35784;
    wire N__35783;
    wire N__35782;
    wire N__35781;
    wire N__35778;
    wire N__35777;
    wire N__35776;
    wire N__35775;
    wire N__35774;
    wire N__35773;
    wire N__35772;
    wire N__35771;
    wire N__35770;
    wire N__35769;
    wire N__35766;
    wire N__35765;
    wire N__35764;
    wire N__35763;
    wire N__35760;
    wire N__35759;
    wire N__35758;
    wire N__35757;
    wire N__35756;
    wire N__35755;
    wire N__35754;
    wire N__35753;
    wire N__35752;
    wire N__35749;
    wire N__35748;
    wire N__35747;
    wire N__35744;
    wire N__35743;
    wire N__35742;
    wire N__35741;
    wire N__35740;
    wire N__35739;
    wire N__35738;
    wire N__35737;
    wire N__35736;
    wire N__35735;
    wire N__35734;
    wire N__35733;
    wire N__35730;
    wire N__35729;
    wire N__35728;
    wire N__35727;
    wire N__35726;
    wire N__35725;
    wire N__35724;
    wire N__35723;
    wire N__35722;
    wire N__35721;
    wire N__35720;
    wire N__35719;
    wire N__35718;
    wire N__35717;
    wire N__35716;
    wire N__35715;
    wire N__35714;
    wire N__35713;
    wire N__35710;
    wire N__35709;
    wire N__35708;
    wire N__35707;
    wire N__35706;
    wire N__35705;
    wire N__35704;
    wire N__35703;
    wire N__35702;
    wire N__35701;
    wire N__35700;
    wire N__35699;
    wire N__35698;
    wire N__35697;
    wire N__35696;
    wire N__35695;
    wire N__35694;
    wire N__35693;
    wire N__35692;
    wire N__35691;
    wire N__35690;
    wire N__35689;
    wire N__35686;
    wire N__35685;
    wire N__35684;
    wire N__35683;
    wire N__35682;
    wire N__35681;
    wire N__35680;
    wire N__35679;
    wire N__35678;
    wire N__35677;
    wire N__35676;
    wire N__35469;
    wire N__35466;
    wire N__35463;
    wire N__35460;
    wire N__35457;
    wire N__35456;
    wire N__35455;
    wire N__35452;
    wire N__35449;
    wire N__35446;
    wire N__35439;
    wire N__35436;
    wire N__35433;
    wire N__35430;
    wire N__35427;
    wire N__35426;
    wire N__35423;
    wire N__35422;
    wire N__35419;
    wire N__35416;
    wire N__35413;
    wire N__35406;
    wire N__35403;
    wire N__35400;
    wire N__35399;
    wire N__35396;
    wire N__35395;
    wire N__35392;
    wire N__35389;
    wire N__35386;
    wire N__35379;
    wire N__35376;
    wire N__35373;
    wire N__35372;
    wire N__35371;
    wire N__35370;
    wire N__35369;
    wire N__35368;
    wire N__35365;
    wire N__35362;
    wire N__35359;
    wire N__35354;
    wire N__35351;
    wire N__35348;
    wire N__35337;
    wire N__35334;
    wire N__35333;
    wire N__35330;
    wire N__35329;
    wire N__35326;
    wire N__35321;
    wire N__35316;
    wire N__35315;
    wire N__35314;
    wire N__35313;
    wire N__35312;
    wire N__35311;
    wire N__35310;
    wire N__35309;
    wire N__35308;
    wire N__35307;
    wire N__35306;
    wire N__35305;
    wire N__35304;
    wire N__35303;
    wire N__35302;
    wire N__35301;
    wire N__35300;
    wire N__35299;
    wire N__35298;
    wire N__35297;
    wire N__35296;
    wire N__35295;
    wire N__35294;
    wire N__35293;
    wire N__35244;
    wire N__35241;
    wire N__35238;
    wire N__35237;
    wire N__35234;
    wire N__35233;
    wire N__35230;
    wire N__35227;
    wire N__35224;
    wire N__35219;
    wire N__35214;
    wire N__35211;
    wire N__35208;
    wire N__35207;
    wire N__35206;
    wire N__35203;
    wire N__35200;
    wire N__35197;
    wire N__35194;
    wire N__35187;
    wire N__35184;
    wire N__35181;
    wire N__35180;
    wire N__35179;
    wire N__35174;
    wire N__35171;
    wire N__35168;
    wire N__35163;
    wire N__35160;
    wire N__35157;
    wire N__35154;
    wire N__35153;
    wire N__35152;
    wire N__35149;
    wire N__35146;
    wire N__35143;
    wire N__35138;
    wire N__35133;
    wire N__35130;
    wire N__35129;
    wire N__35128;
    wire N__35125;
    wire N__35122;
    wire N__35119;
    wire N__35112;
    wire N__35109;
    wire N__35108;
    wire N__35107;
    wire N__35104;
    wire N__35101;
    wire N__35096;
    wire N__35091;
    wire N__35088;
    wire N__35087;
    wire N__35086;
    wire N__35085;
    wire N__35076;
    wire N__35073;
    wire N__35070;
    wire N__35067;
    wire N__35064;
    wire N__35061;
    wire N__35060;
    wire N__35057;
    wire N__35054;
    wire N__35051;
    wire N__35050;
    wire N__35047;
    wire N__35044;
    wire N__35041;
    wire N__35038;
    wire N__35033;
    wire N__35030;
    wire N__35025;
    wire N__35024;
    wire N__35021;
    wire N__35018;
    wire N__35015;
    wire N__35012;
    wire N__35009;
    wire N__35008;
    wire N__35005;
    wire N__35002;
    wire N__34999;
    wire N__34994;
    wire N__34989;
    wire N__34986;
    wire N__34983;
    wire N__34980;
    wire N__34979;
    wire N__34978;
    wire N__34975;
    wire N__34972;
    wire N__34969;
    wire N__34966;
    wire N__34961;
    wire N__34958;
    wire N__34953;
    wire N__34950;
    wire N__34947;
    wire N__34944;
    wire N__34941;
    wire N__34938;
    wire N__34935;
    wire N__34932;
    wire N__34929;
    wire N__34926;
    wire N__34923;
    wire N__34920;
    wire N__34917;
    wire N__34914;
    wire N__34911;
    wire N__34908;
    wire N__34905;
    wire N__34902;
    wire N__34899;
    wire N__34896;
    wire N__34895;
    wire N__34894;
    wire N__34893;
    wire N__34890;
    wire N__34889;
    wire N__34886;
    wire N__34885;
    wire N__34884;
    wire N__34883;
    wire N__34880;
    wire N__34877;
    wire N__34874;
    wire N__34871;
    wire N__34870;
    wire N__34867;
    wire N__34864;
    wire N__34863;
    wire N__34862;
    wire N__34859;
    wire N__34856;
    wire N__34851;
    wire N__34848;
    wire N__34845;
    wire N__34842;
    wire N__34839;
    wire N__34836;
    wire N__34833;
    wire N__34828;
    wire N__34823;
    wire N__34818;
    wire N__34803;
    wire N__34802;
    wire N__34799;
    wire N__34796;
    wire N__34793;
    wire N__34790;
    wire N__34789;
    wire N__34784;
    wire N__34781;
    wire N__34778;
    wire N__34773;
    wire N__34772;
    wire N__34771;
    wire N__34768;
    wire N__34765;
    wire N__34764;
    wire N__34763;
    wire N__34762;
    wire N__34761;
    wire N__34758;
    wire N__34755;
    wire N__34752;
    wire N__34749;
    wire N__34746;
    wire N__34743;
    wire N__34742;
    wire N__34739;
    wire N__34734;
    wire N__34733;
    wire N__34732;
    wire N__34731;
    wire N__34728;
    wire N__34725;
    wire N__34722;
    wire N__34719;
    wire N__34716;
    wire N__34711;
    wire N__34706;
    wire N__34703;
    wire N__34696;
    wire N__34683;
    wire N__34680;
    wire N__34677;
    wire N__34676;
    wire N__34675;
    wire N__34672;
    wire N__34669;
    wire N__34666;
    wire N__34663;
    wire N__34660;
    wire N__34655;
    wire N__34650;
    wire N__34649;
    wire N__34646;
    wire N__34645;
    wire N__34642;
    wire N__34639;
    wire N__34636;
    wire N__34633;
    wire N__34628;
    wire N__34625;
    wire N__34622;
    wire N__34619;
    wire N__34614;
    wire N__34611;
    wire N__34610;
    wire N__34609;
    wire N__34606;
    wire N__34603;
    wire N__34600;
    wire N__34597;
    wire N__34594;
    wire N__34591;
    wire N__34588;
    wire N__34581;
    wire N__34578;
    wire N__34575;
    wire N__34572;
    wire N__34571;
    wire N__34568;
    wire N__34567;
    wire N__34564;
    wire N__34561;
    wire N__34558;
    wire N__34551;
    wire N__34550;
    wire N__34549;
    wire N__34546;
    wire N__34541;
    wire N__34536;
    wire N__34535;
    wire N__34534;
    wire N__34531;
    wire N__34528;
    wire N__34525;
    wire N__34520;
    wire N__34515;
    wire N__34512;
    wire N__34511;
    wire N__34508;
    wire N__34505;
    wire N__34502;
    wire N__34501;
    wire N__34500;
    wire N__34497;
    wire N__34496;
    wire N__34495;
    wire N__34492;
    wire N__34489;
    wire N__34486;
    wire N__34483;
    wire N__34480;
    wire N__34477;
    wire N__34472;
    wire N__34471;
    wire N__34470;
    wire N__34469;
    wire N__34466;
    wire N__34459;
    wire N__34456;
    wire N__34453;
    wire N__34450;
    wire N__34447;
    wire N__34442;
    wire N__34439;
    wire N__34432;
    wire N__34429;
    wire N__34426;
    wire N__34423;
    wire N__34416;
    wire N__34415;
    wire N__34414;
    wire N__34413;
    wire N__34410;
    wire N__34407;
    wire N__34404;
    wire N__34403;
    wire N__34402;
    wire N__34401;
    wire N__34400;
    wire N__34399;
    wire N__34396;
    wire N__34395;
    wire N__34394;
    wire N__34391;
    wire N__34388;
    wire N__34385;
    wire N__34382;
    wire N__34379;
    wire N__34378;
    wire N__34375;
    wire N__34374;
    wire N__34373;
    wire N__34370;
    wire N__34367;
    wire N__34366;
    wire N__34365;
    wire N__34362;
    wire N__34359;
    wire N__34356;
    wire N__34351;
    wire N__34346;
    wire N__34343;
    wire N__34340;
    wire N__34337;
    wire N__34332;
    wire N__34329;
    wire N__34326;
    wire N__34323;
    wire N__34320;
    wire N__34317;
    wire N__34312;
    wire N__34309;
    wire N__34304;
    wire N__34301;
    wire N__34298;
    wire N__34295;
    wire N__34292;
    wire N__34285;
    wire N__34276;
    wire N__34269;
    wire N__34264;
    wire N__34257;
    wire N__34254;
    wire N__34251;
    wire N__34250;
    wire N__34249;
    wire N__34246;
    wire N__34243;
    wire N__34240;
    wire N__34237;
    wire N__34234;
    wire N__34229;
    wire N__34224;
    wire N__34221;
    wire N__34218;
    wire N__34217;
    wire N__34214;
    wire N__34211;
    wire N__34208;
    wire N__34207;
    wire N__34204;
    wire N__34201;
    wire N__34198;
    wire N__34195;
    wire N__34192;
    wire N__34189;
    wire N__34186;
    wire N__34183;
    wire N__34176;
    wire N__34173;
    wire N__34170;
    wire N__34167;
    wire N__34164;
    wire N__34163;
    wire N__34160;
    wire N__34157;
    wire N__34154;
    wire N__34153;
    wire N__34150;
    wire N__34147;
    wire N__34144;
    wire N__34141;
    wire N__34134;
    wire N__34131;
    wire N__34128;
    wire N__34125;
    wire N__34122;
    wire N__34121;
    wire N__34118;
    wire N__34115;
    wire N__34114;
    wire N__34111;
    wire N__34108;
    wire N__34105;
    wire N__34098;
    wire N__34095;
    wire N__34092;
    wire N__34089;
    wire N__34088;
    wire N__34087;
    wire N__34086;
    wire N__34085;
    wire N__34082;
    wire N__34081;
    wire N__34078;
    wire N__34077;
    wire N__34074;
    wire N__34071;
    wire N__34068;
    wire N__34065;
    wire N__34062;
    wire N__34061;
    wire N__34054;
    wire N__34049;
    wire N__34048;
    wire N__34047;
    wire N__34046;
    wire N__34043;
    wire N__34038;
    wire N__34033;
    wire N__34032;
    wire N__34031;
    wire N__34030;
    wire N__34029;
    wire N__34028;
    wire N__34025;
    wire N__34022;
    wire N__34019;
    wire N__34014;
    wire N__34011;
    wire N__34002;
    wire N__33997;
    wire N__33984;
    wire N__33981;
    wire N__33980;
    wire N__33977;
    wire N__33974;
    wire N__33971;
    wire N__33970;
    wire N__33967;
    wire N__33964;
    wire N__33961;
    wire N__33958;
    wire N__33951;
    wire N__33950;
    wire N__33949;
    wire N__33946;
    wire N__33945;
    wire N__33944;
    wire N__33943;
    wire N__33942;
    wire N__33939;
    wire N__33932;
    wire N__33927;
    wire N__33926;
    wire N__33925;
    wire N__33924;
    wire N__33919;
    wire N__33914;
    wire N__33913;
    wire N__33910;
    wire N__33909;
    wire N__33906;
    wire N__33905;
    wire N__33904;
    wire N__33903;
    wire N__33900;
    wire N__33897;
    wire N__33894;
    wire N__33883;
    wire N__33878;
    wire N__33867;
    wire N__33864;
    wire N__33861;
    wire N__33858;
    wire N__33857;
    wire N__33856;
    wire N__33855;
    wire N__33852;
    wire N__33851;
    wire N__33850;
    wire N__33849;
    wire N__33848;
    wire N__33847;
    wire N__33846;
    wire N__33843;
    wire N__33842;
    wire N__33837;
    wire N__33834;
    wire N__33831;
    wire N__33830;
    wire N__33829;
    wire N__33828;
    wire N__33827;
    wire N__33826;
    wire N__33823;
    wire N__33822;
    wire N__33819;
    wire N__33816;
    wire N__33813;
    wire N__33810;
    wire N__33807;
    wire N__33804;
    wire N__33801;
    wire N__33796;
    wire N__33793;
    wire N__33788;
    wire N__33785;
    wire N__33784;
    wire N__33783;
    wire N__33780;
    wire N__33777;
    wire N__33774;
    wire N__33771;
    wire N__33762;
    wire N__33761;
    wire N__33760;
    wire N__33759;
    wire N__33752;
    wire N__33751;
    wire N__33750;
    wire N__33749;
    wire N__33744;
    wire N__33741;
    wire N__33736;
    wire N__33733;
    wire N__33730;
    wire N__33723;
    wire N__33716;
    wire N__33713;
    wire N__33708;
    wire N__33705;
    wire N__33702;
    wire N__33699;
    wire N__33690;
    wire N__33685;
    wire N__33672;
    wire N__33671;
    wire N__33670;
    wire N__33667;
    wire N__33666;
    wire N__33663;
    wire N__33662;
    wire N__33661;
    wire N__33660;
    wire N__33659;
    wire N__33658;
    wire N__33657;
    wire N__33656;
    wire N__33653;
    wire N__33652;
    wire N__33651;
    wire N__33648;
    wire N__33645;
    wire N__33640;
    wire N__33639;
    wire N__33638;
    wire N__33637;
    wire N__33634;
    wire N__33631;
    wire N__33628;
    wire N__33623;
    wire N__33620;
    wire N__33619;
    wire N__33616;
    wire N__33611;
    wire N__33604;
    wire N__33601;
    wire N__33600;
    wire N__33599;
    wire N__33596;
    wire N__33593;
    wire N__33590;
    wire N__33587;
    wire N__33586;
    wire N__33583;
    wire N__33578;
    wire N__33575;
    wire N__33572;
    wire N__33565;
    wire N__33562;
    wire N__33561;
    wire N__33560;
    wire N__33559;
    wire N__33558;
    wire N__33557;
    wire N__33554;
    wire N__33549;
    wire N__33546;
    wire N__33543;
    wire N__33540;
    wire N__33537;
    wire N__33534;
    wire N__33531;
    wire N__33526;
    wire N__33521;
    wire N__33518;
    wire N__33511;
    wire N__33508;
    wire N__33503;
    wire N__33500;
    wire N__33493;
    wire N__33490;
    wire N__33487;
    wire N__33468;
    wire N__33467;
    wire N__33466;
    wire N__33465;
    wire N__33464;
    wire N__33463;
    wire N__33460;
    wire N__33459;
    wire N__33458;
    wire N__33457;
    wire N__33456;
    wire N__33453;
    wire N__33452;
    wire N__33451;
    wire N__33450;
    wire N__33449;
    wire N__33448;
    wire N__33447;
    wire N__33446;
    wire N__33443;
    wire N__33442;
    wire N__33441;
    wire N__33440;
    wire N__33437;
    wire N__33436;
    wire N__33433;
    wire N__33432;
    wire N__33429;
    wire N__33426;
    wire N__33421;
    wire N__33416;
    wire N__33413;
    wire N__33410;
    wire N__33407;
    wire N__33404;
    wire N__33401;
    wire N__33400;
    wire N__33397;
    wire N__33394;
    wire N__33391;
    wire N__33388;
    wire N__33385;
    wire N__33382;
    wire N__33377;
    wire N__33374;
    wire N__33371;
    wire N__33368;
    wire N__33367;
    wire N__33364;
    wire N__33357;
    wire N__33354;
    wire N__33351;
    wire N__33346;
    wire N__33343;
    wire N__33340;
    wire N__33337;
    wire N__33332;
    wire N__33329;
    wire N__33326;
    wire N__33323;
    wire N__33316;
    wire N__33311;
    wire N__33304;
    wire N__33301;
    wire N__33298;
    wire N__33295;
    wire N__33292;
    wire N__33287;
    wire N__33284;
    wire N__33283;
    wire N__33276;
    wire N__33267;
    wire N__33264;
    wire N__33259;
    wire N__33256;
    wire N__33253;
    wire N__33246;
    wire N__33241;
    wire N__33234;
    wire N__33233;
    wire N__33232;
    wire N__33231;
    wire N__33226;
    wire N__33225;
    wire N__33224;
    wire N__33221;
    wire N__33218;
    wire N__33215;
    wire N__33214;
    wire N__33211;
    wire N__33208;
    wire N__33207;
    wire N__33204;
    wire N__33203;
    wire N__33200;
    wire N__33197;
    wire N__33194;
    wire N__33193;
    wire N__33192;
    wire N__33189;
    wire N__33186;
    wire N__33183;
    wire N__33180;
    wire N__33177;
    wire N__33174;
    wire N__33169;
    wire N__33164;
    wire N__33157;
    wire N__33154;
    wire N__33151;
    wire N__33144;
    wire N__33141;
    wire N__33132;
    wire N__33131;
    wire N__33130;
    wire N__33129;
    wire N__33128;
    wire N__33127;
    wire N__33126;
    wire N__33121;
    wire N__33120;
    wire N__33117;
    wire N__33116;
    wire N__33115;
    wire N__33114;
    wire N__33113;
    wire N__33112;
    wire N__33111;
    wire N__33110;
    wire N__33109;
    wire N__33104;
    wire N__33103;
    wire N__33102;
    wire N__33101;
    wire N__33100;
    wire N__33097;
    wire N__33094;
    wire N__33091;
    wire N__33088;
    wire N__33085;
    wire N__33074;
    wire N__33069;
    wire N__33066;
    wire N__33063;
    wire N__33054;
    wire N__33053;
    wire N__33052;
    wire N__33049;
    wire N__33048;
    wire N__33047;
    wire N__33046;
    wire N__33045;
    wire N__33044;
    wire N__33039;
    wire N__33030;
    wire N__33027;
    wire N__33022;
    wire N__33019;
    wire N__33016;
    wire N__33015;
    wire N__33014;
    wire N__33013;
    wire N__33012;
    wire N__33009;
    wire N__33000;
    wire N__32997;
    wire N__32992;
    wire N__32987;
    wire N__32974;
    wire N__32969;
    wire N__32958;
    wire N__32955;
    wire N__32952;
    wire N__32949;
    wire N__32948;
    wire N__32947;
    wire N__32946;
    wire N__32945;
    wire N__32944;
    wire N__32941;
    wire N__32938;
    wire N__32935;
    wire N__32930;
    wire N__32927;
    wire N__32926;
    wire N__32923;
    wire N__32922;
    wire N__32919;
    wire N__32916;
    wire N__32911;
    wire N__32910;
    wire N__32909;
    wire N__32908;
    wire N__32905;
    wire N__32902;
    wire N__32899;
    wire N__32892;
    wire N__32887;
    wire N__32884;
    wire N__32871;
    wire N__32868;
    wire N__32867;
    wire N__32866;
    wire N__32863;
    wire N__32860;
    wire N__32857;
    wire N__32854;
    wire N__32851;
    wire N__32848;
    wire N__32841;
    wire N__32840;
    wire N__32839;
    wire N__32836;
    wire N__32835;
    wire N__32832;
    wire N__32831;
    wire N__32830;
    wire N__32827;
    wire N__32822;
    wire N__32819;
    wire N__32818;
    wire N__32815;
    wire N__32812;
    wire N__32811;
    wire N__32810;
    wire N__32807;
    wire N__32802;
    wire N__32801;
    wire N__32800;
    wire N__32797;
    wire N__32794;
    wire N__32791;
    wire N__32788;
    wire N__32785;
    wire N__32780;
    wire N__32775;
    wire N__32772;
    wire N__32757;
    wire N__32754;
    wire N__32751;
    wire N__32750;
    wire N__32747;
    wire N__32744;
    wire N__32739;
    wire N__32736;
    wire N__32733;
    wire N__32730;
    wire N__32729;
    wire N__32726;
    wire N__32723;
    wire N__32720;
    wire N__32717;
    wire N__32716;
    wire N__32713;
    wire N__32710;
    wire N__32707;
    wire N__32700;
    wire N__32697;
    wire N__32694;
    wire N__32691;
    wire N__32688;
    wire N__32687;
    wire N__32684;
    wire N__32683;
    wire N__32680;
    wire N__32675;
    wire N__32670;
    wire N__32667;
    wire N__32664;
    wire N__32661;
    wire N__32658;
    wire N__32657;
    wire N__32654;
    wire N__32651;
    wire N__32650;
    wire N__32645;
    wire N__32642;
    wire N__32637;
    wire N__32634;
    wire N__32631;
    wire N__32628;
    wire N__32627;
    wire N__32622;
    wire N__32619;
    wire N__32616;
    wire N__32613;
    wire N__32610;
    wire N__32607;
    wire N__32604;
    wire N__32601;
    wire N__32598;
    wire N__32595;
    wire N__32592;
    wire N__32591;
    wire N__32590;
    wire N__32589;
    wire N__32588;
    wire N__32587;
    wire N__32586;
    wire N__32585;
    wire N__32584;
    wire N__32583;
    wire N__32582;
    wire N__32581;
    wire N__32580;
    wire N__32579;
    wire N__32578;
    wire N__32577;
    wire N__32576;
    wire N__32575;
    wire N__32574;
    wire N__32573;
    wire N__32572;
    wire N__32571;
    wire N__32570;
    wire N__32569;
    wire N__32568;
    wire N__32567;
    wire N__32566;
    wire N__32563;
    wire N__32560;
    wire N__32557;
    wire N__32554;
    wire N__32551;
    wire N__32548;
    wire N__32545;
    wire N__32544;
    wire N__32543;
    wire N__32542;
    wire N__32541;
    wire N__32540;
    wire N__32539;
    wire N__32538;
    wire N__32535;
    wire N__32534;
    wire N__32531;
    wire N__32528;
    wire N__32525;
    wire N__32522;
    wire N__32519;
    wire N__32518;
    wire N__32515;
    wire N__32512;
    wire N__32509;
    wire N__32506;
    wire N__32503;
    wire N__32500;
    wire N__32497;
    wire N__32496;
    wire N__32495;
    wire N__32494;
    wire N__32491;
    wire N__32488;
    wire N__32485;
    wire N__32482;
    wire N__32479;
    wire N__32476;
    wire N__32473;
    wire N__32472;
    wire N__32471;
    wire N__32470;
    wire N__32469;
    wire N__32468;
    wire N__32467;
    wire N__32466;
    wire N__32457;
    wire N__32450;
    wire N__32447;
    wire N__32444;
    wire N__32441;
    wire N__32438;
    wire N__32435;
    wire N__32432;
    wire N__32429;
    wire N__32418;
    wire N__32413;
    wire N__32412;
    wire N__32411;
    wire N__32410;
    wire N__32407;
    wire N__32398;
    wire N__32391;
    wire N__32390;
    wire N__32387;
    wire N__32384;
    wire N__32383;
    wire N__32382;
    wire N__32379;
    wire N__32370;
    wire N__32363;
    wire N__32360;
    wire N__32357;
    wire N__32354;
    wire N__32351;
    wire N__32348;
    wire N__32345;
    wire N__32342;
    wire N__32339;
    wire N__32336;
    wire N__32327;
    wire N__32320;
    wire N__32315;
    wire N__32314;
    wire N__32311;
    wire N__32308;
    wire N__32307;
    wire N__32306;
    wire N__32305;
    wire N__32302;
    wire N__32299;
    wire N__32294;
    wire N__32281;
    wire N__32276;
    wire N__32267;
    wire N__32260;
    wire N__32255;
    wire N__32250;
    wire N__32247;
    wire N__32232;
    wire N__32229;
    wire N__32224;
    wire N__32221;
    wire N__32216;
    wire N__32211;
    wire N__32208;
    wire N__32205;
    wire N__32202;
    wire N__32199;
    wire N__32194;
    wire N__32191;
    wire N__32186;
    wire N__32179;
    wire N__32172;
    wire N__32169;
    wire N__32166;
    wire N__32163;
    wire N__32160;
    wire N__32157;
    wire N__32154;
    wire N__32151;
    wire N__32148;
    wire N__32145;
    wire N__32142;
    wire N__32141;
    wire N__32138;
    wire N__32135;
    wire N__32130;
    wire N__32127;
    wire N__32124;
    wire N__32121;
    wire N__32118;
    wire N__32115;
    wire N__32112;
    wire N__32109;
    wire N__32106;
    wire N__32103;
    wire N__32100;
    wire N__32097;
    wire N__32094;
    wire N__32091;
    wire N__32088;
    wire N__32087;
    wire N__32086;
    wire N__32085;
    wire N__32084;
    wire N__32083;
    wire N__32082;
    wire N__32079;
    wire N__32074;
    wire N__32073;
    wire N__32072;
    wire N__32069;
    wire N__32066;
    wire N__32063;
    wire N__32060;
    wire N__32057;
    wire N__32054;
    wire N__32051;
    wire N__32050;
    wire N__32047;
    wire N__32044;
    wire N__32043;
    wire N__32040;
    wire N__32037;
    wire N__32034;
    wire N__32033;
    wire N__32026;
    wire N__32023;
    wire N__32022;
    wire N__32021;
    wire N__32020;
    wire N__32017;
    wire N__32014;
    wire N__32011;
    wire N__32008;
    wire N__32005;
    wire N__32002;
    wire N__31999;
    wire N__31994;
    wire N__31989;
    wire N__31986;
    wire N__31985;
    wire N__31978;
    wire N__31973;
    wire N__31970;
    wire N__31967;
    wire N__31964;
    wire N__31959;
    wire N__31956;
    wire N__31951;
    wire N__31942;
    wire N__31935;
    wire N__31932;
    wire N__31929;
    wire N__31926;
    wire N__31923;
    wire N__31920;
    wire N__31919;
    wire N__31918;
    wire N__31917;
    wire N__31916;
    wire N__31913;
    wire N__31910;
    wire N__31909;
    wire N__31908;
    wire N__31905;
    wire N__31904;
    wire N__31903;
    wire N__31900;
    wire N__31897;
    wire N__31896;
    wire N__31895;
    wire N__31894;
    wire N__31891;
    wire N__31888;
    wire N__31885;
    wire N__31882;
    wire N__31879;
    wire N__31878;
    wire N__31875;
    wire N__31872;
    wire N__31871;
    wire N__31868;
    wire N__31865;
    wire N__31862;
    wire N__31859;
    wire N__31858;
    wire N__31857;
    wire N__31854;
    wire N__31849;
    wire N__31846;
    wire N__31843;
    wire N__31840;
    wire N__31837;
    wire N__31832;
    wire N__31829;
    wire N__31826;
    wire N__31823;
    wire N__31820;
    wire N__31817;
    wire N__31814;
    wire N__31811;
    wire N__31808;
    wire N__31801;
    wire N__31798;
    wire N__31795;
    wire N__31792;
    wire N__31789;
    wire N__31786;
    wire N__31779;
    wire N__31776;
    wire N__31773;
    wire N__31768;
    wire N__31765;
    wire N__31758;
    wire N__31753;
    wire N__31746;
    wire N__31737;
    wire N__31734;
    wire N__31731;
    wire N__31728;
    wire N__31725;
    wire N__31722;
    wire N__31719;
    wire N__31716;
    wire N__31713;
    wire N__31710;
    wire N__31707;
    wire N__31704;
    wire N__31701;
    wire N__31698;
    wire N__31695;
    wire N__31692;
    wire N__31691;
    wire N__31690;
    wire N__31683;
    wire N__31680;
    wire N__31677;
    wire N__31676;
    wire N__31671;
    wire N__31668;
    wire N__31665;
    wire N__31664;
    wire N__31661;
    wire N__31658;
    wire N__31657;
    wire N__31656;
    wire N__31647;
    wire N__31644;
    wire N__31643;
    wire N__31642;
    wire N__31641;
    wire N__31632;
    wire N__31629;
    wire N__31626;
    wire N__31623;
    wire N__31620;
    wire N__31617;
    wire N__31614;
    wire N__31611;
    wire N__31608;
    wire N__31605;
    wire N__31604;
    wire N__31603;
    wire N__31600;
    wire N__31597;
    wire N__31594;
    wire N__31593;
    wire N__31592;
    wire N__31591;
    wire N__31590;
    wire N__31589;
    wire N__31588;
    wire N__31587;
    wire N__31586;
    wire N__31585;
    wire N__31584;
    wire N__31583;
    wire N__31580;
    wire N__31577;
    wire N__31574;
    wire N__31571;
    wire N__31568;
    wire N__31565;
    wire N__31560;
    wire N__31555;
    wire N__31550;
    wire N__31547;
    wire N__31544;
    wire N__31543;
    wire N__31542;
    wire N__31539;
    wire N__31534;
    wire N__31531;
    wire N__31528;
    wire N__31525;
    wire N__31520;
    wire N__31517;
    wire N__31512;
    wire N__31509;
    wire N__31506;
    wire N__31501;
    wire N__31498;
    wire N__31493;
    wire N__31488;
    wire N__31483;
    wire N__31480;
    wire N__31477;
    wire N__31474;
    wire N__31469;
    wire N__31464;
    wire N__31455;
    wire N__31452;
    wire N__31449;
    wire N__31446;
    wire N__31443;
    wire N__31440;
    wire N__31439;
    wire N__31438;
    wire N__31437;
    wire N__31436;
    wire N__31435;
    wire N__31434;
    wire N__31431;
    wire N__31430;
    wire N__31429;
    wire N__31426;
    wire N__31423;
    wire N__31422;
    wire N__31419;
    wire N__31416;
    wire N__31413;
    wire N__31412;
    wire N__31411;
    wire N__31408;
    wire N__31407;
    wire N__31404;
    wire N__31395;
    wire N__31392;
    wire N__31389;
    wire N__31386;
    wire N__31383;
    wire N__31382;
    wire N__31379;
    wire N__31378;
    wire N__31375;
    wire N__31374;
    wire N__31369;
    wire N__31364;
    wire N__31361;
    wire N__31358;
    wire N__31355;
    wire N__31352;
    wire N__31349;
    wire N__31346;
    wire N__31343;
    wire N__31340;
    wire N__31337;
    wire N__31332;
    wire N__31325;
    wire N__31322;
    wire N__31317;
    wire N__31314;
    wire N__31311;
    wire N__31308;
    wire N__31303;
    wire N__31298;
    wire N__31287;
    wire N__31284;
    wire N__31281;
    wire N__31280;
    wire N__31279;
    wire N__31278;
    wire N__31275;
    wire N__31272;
    wire N__31271;
    wire N__31268;
    wire N__31265;
    wire N__31264;
    wire N__31261;
    wire N__31258;
    wire N__31257;
    wire N__31256;
    wire N__31253;
    wire N__31252;
    wire N__31249;
    wire N__31248;
    wire N__31247;
    wire N__31244;
    wire N__31241;
    wire N__31240;
    wire N__31239;
    wire N__31236;
    wire N__31233;
    wire N__31230;
    wire N__31227;
    wire N__31224;
    wire N__31221;
    wire N__31220;
    wire N__31219;
    wire N__31218;
    wire N__31215;
    wire N__31212;
    wire N__31209;
    wire N__31206;
    wire N__31203;
    wire N__31200;
    wire N__31197;
    wire N__31190;
    wire N__31187;
    wire N__31182;
    wire N__31175;
    wire N__31168;
    wire N__31163;
    wire N__31158;
    wire N__31153;
    wire N__31146;
    wire N__31137;
    wire N__31134;
    wire N__31131;
    wire N__31128;
    wire N__31125;
    wire N__31124;
    wire N__31121;
    wire N__31120;
    wire N__31119;
    wire N__31118;
    wire N__31115;
    wire N__31114;
    wire N__31113;
    wire N__31112;
    wire N__31111;
    wire N__31110;
    wire N__31109;
    wire N__31108;
    wire N__31107;
    wire N__31104;
    wire N__31101;
    wire N__31098;
    wire N__31095;
    wire N__31094;
    wire N__31091;
    wire N__31088;
    wire N__31087;
    wire N__31082;
    wire N__31079;
    wire N__31076;
    wire N__31073;
    wire N__31070;
    wire N__31067;
    wire N__31064;
    wire N__31063;
    wire N__31060;
    wire N__31057;
    wire N__31054;
    wire N__31051;
    wire N__31048;
    wire N__31045;
    wire N__31042;
    wire N__31037;
    wire N__31032;
    wire N__31027;
    wire N__31024;
    wire N__31021;
    wire N__31018;
    wire N__31011;
    wire N__31004;
    wire N__31001;
    wire N__30996;
    wire N__30991;
    wire N__30988;
    wire N__30981;
    wire N__30978;
    wire N__30969;
    wire N__30966;
    wire N__30963;
    wire N__30960;
    wire N__30957;
    wire N__30954;
    wire N__30951;
    wire N__30948;
    wire N__30947;
    wire N__30944;
    wire N__30943;
    wire N__30940;
    wire N__30937;
    wire N__30934;
    wire N__30931;
    wire N__30928;
    wire N__30925;
    wire N__30918;
    wire N__30915;
    wire N__30912;
    wire N__30909;
    wire N__30908;
    wire N__30907;
    wire N__30904;
    wire N__30901;
    wire N__30898;
    wire N__30895;
    wire N__30892;
    wire N__30885;
    wire N__30882;
    wire N__30879;
    wire N__30878;
    wire N__30877;
    wire N__30874;
    wire N__30871;
    wire N__30868;
    wire N__30865;
    wire N__30862;
    wire N__30857;
    wire N__30854;
    wire N__30849;
    wire N__30846;
    wire N__30845;
    wire N__30842;
    wire N__30839;
    wire N__30838;
    wire N__30835;
    wire N__30832;
    wire N__30829;
    wire N__30826;
    wire N__30823;
    wire N__30818;
    wire N__30815;
    wire N__30810;
    wire N__30809;
    wire N__30806;
    wire N__30803;
    wire N__30800;
    wire N__30799;
    wire N__30796;
    wire N__30793;
    wire N__30790;
    wire N__30785;
    wire N__30780;
    wire N__30777;
    wire N__30776;
    wire N__30773;
    wire N__30770;
    wire N__30769;
    wire N__30766;
    wire N__30763;
    wire N__30760;
    wire N__30757;
    wire N__30754;
    wire N__30747;
    wire N__30744;
    wire N__30741;
    wire N__30738;
    wire N__30735;
    wire N__30732;
    wire N__30729;
    wire N__30726;
    wire N__30723;
    wire N__30720;
    wire N__30717;
    wire N__30714;
    wire N__30711;
    wire N__30710;
    wire N__30707;
    wire N__30704;
    wire N__30703;
    wire N__30700;
    wire N__30697;
    wire N__30694;
    wire N__30691;
    wire N__30688;
    wire N__30685;
    wire N__30680;
    wire N__30675;
    wire N__30672;
    wire N__30669;
    wire N__30668;
    wire N__30665;
    wire N__30662;
    wire N__30661;
    wire N__30658;
    wire N__30655;
    wire N__30652;
    wire N__30649;
    wire N__30642;
    wire N__30639;
    wire N__30638;
    wire N__30635;
    wire N__30634;
    wire N__30631;
    wire N__30628;
    wire N__30625;
    wire N__30622;
    wire N__30621;
    wire N__30616;
    wire N__30613;
    wire N__30610;
    wire N__30607;
    wire N__30600;
    wire N__30597;
    wire N__30594;
    wire N__30591;
    wire N__30588;
    wire N__30585;
    wire N__30582;
    wire N__30581;
    wire N__30576;
    wire N__30573;
    wire N__30570;
    wire N__30569;
    wire N__30568;
    wire N__30565;
    wire N__30562;
    wire N__30559;
    wire N__30556;
    wire N__30551;
    wire N__30548;
    wire N__30545;
    wire N__30542;
    wire N__30539;
    wire N__30534;
    wire N__30531;
    wire N__30530;
    wire N__30527;
    wire N__30526;
    wire N__30523;
    wire N__30520;
    wire N__30517;
    wire N__30514;
    wire N__30511;
    wire N__30508;
    wire N__30505;
    wire N__30502;
    wire N__30499;
    wire N__30492;
    wire N__30489;
    wire N__30486;
    wire N__30483;
    wire N__30480;
    wire N__30477;
    wire N__30474;
    wire N__30471;
    wire N__30468;
    wire N__30465;
    wire N__30462;
    wire N__30461;
    wire N__30460;
    wire N__30457;
    wire N__30454;
    wire N__30451;
    wire N__30446;
    wire N__30443;
    wire N__30440;
    wire N__30437;
    wire N__30434;
    wire N__30431;
    wire N__30426;
    wire N__30423;
    wire N__30422;
    wire N__30419;
    wire N__30418;
    wire N__30415;
    wire N__30412;
    wire N__30409;
    wire N__30406;
    wire N__30403;
    wire N__30400;
    wire N__30397;
    wire N__30392;
    wire N__30387;
    wire N__30386;
    wire N__30383;
    wire N__30380;
    wire N__30379;
    wire N__30376;
    wire N__30373;
    wire N__30370;
    wire N__30367;
    wire N__30362;
    wire N__30357;
    wire N__30354;
    wire N__30353;
    wire N__30350;
    wire N__30347;
    wire N__30346;
    wire N__30341;
    wire N__30338;
    wire N__30335;
    wire N__30332;
    wire N__30327;
    wire N__30324;
    wire N__30321;
    wire N__30318;
    wire N__30317;
    wire N__30314;
    wire N__30311;
    wire N__30308;
    wire N__30305;
    wire N__30300;
    wire N__30299;
    wire N__30296;
    wire N__30293;
    wire N__30290;
    wire N__30285;
    wire N__30284;
    wire N__30281;
    wire N__30278;
    wire N__30275;
    wire N__30272;
    wire N__30269;
    wire N__30268;
    wire N__30265;
    wire N__30262;
    wire N__30259;
    wire N__30256;
    wire N__30253;
    wire N__30248;
    wire N__30243;
    wire N__30240;
    wire N__30237;
    wire N__30234;
    wire N__30231;
    wire N__30228;
    wire N__30227;
    wire N__30226;
    wire N__30223;
    wire N__30218;
    wire N__30213;
    wire N__30210;
    wire N__30207;
    wire N__30204;
    wire N__30201;
    wire N__30198;
    wire N__30195;
    wire N__30194;
    wire N__30193;
    wire N__30190;
    wire N__30185;
    wire N__30180;
    wire N__30177;
    wire N__30174;
    wire N__30171;
    wire N__30168;
    wire N__30165;
    wire N__30162;
    wire N__30161;
    wire N__30158;
    wire N__30157;
    wire N__30154;
    wire N__30151;
    wire N__30148;
    wire N__30145;
    wire N__30140;
    wire N__30137;
    wire N__30134;
    wire N__30129;
    wire N__30126;
    wire N__30123;
    wire N__30120;
    wire N__30117;
    wire N__30114;
    wire N__30111;
    wire N__30108;
    wire N__30105;
    wire N__30102;
    wire N__30099;
    wire N__30098;
    wire N__30097;
    wire N__30094;
    wire N__30091;
    wire N__30088;
    wire N__30083;
    wire N__30080;
    wire N__30075;
    wire N__30072;
    wire N__30069;
    wire N__30066;
    wire N__30063;
    wire N__30060;
    wire N__30057;
    wire N__30054;
    wire N__30053;
    wire N__30050;
    wire N__30049;
    wire N__30046;
    wire N__30043;
    wire N__30040;
    wire N__30033;
    wire N__30030;
    wire N__30027;
    wire N__30024;
    wire N__30021;
    wire N__30018;
    wire N__30015;
    wire N__30014;
    wire N__30013;
    wire N__30010;
    wire N__30007;
    wire N__30002;
    wire N__29997;
    wire N__29994;
    wire N__29991;
    wire N__29988;
    wire N__29985;
    wire N__29982;
    wire N__29979;
    wire N__29976;
    wire N__29973;
    wire N__29970;
    wire N__29969;
    wire N__29966;
    wire N__29965;
    wire N__29962;
    wire N__29959;
    wire N__29956;
    wire N__29953;
    wire N__29950;
    wire N__29947;
    wire N__29944;
    wire N__29941;
    wire N__29934;
    wire N__29931;
    wire N__29928;
    wire N__29925;
    wire N__29922;
    wire N__29919;
    wire N__29916;
    wire N__29913;
    wire N__29910;
    wire N__29907;
    wire N__29906;
    wire N__29903;
    wire N__29900;
    wire N__29897;
    wire N__29892;
    wire N__29889;
    wire N__29886;
    wire N__29883;
    wire N__29880;
    wire N__29877;
    wire N__29874;
    wire N__29871;
    wire N__29868;
    wire N__29865;
    wire N__29862;
    wire N__29859;
    wire N__29856;
    wire N__29853;
    wire N__29850;
    wire N__29847;
    wire N__29844;
    wire N__29841;
    wire N__29838;
    wire N__29835;
    wire N__29832;
    wire N__29829;
    wire N__29826;
    wire N__29823;
    wire N__29820;
    wire N__29817;
    wire N__29814;
    wire N__29811;
    wire N__29808;
    wire N__29805;
    wire N__29802;
    wire N__29799;
    wire N__29796;
    wire N__29793;
    wire N__29790;
    wire N__29787;
    wire N__29784;
    wire N__29781;
    wire N__29778;
    wire N__29775;
    wire N__29772;
    wire N__29771;
    wire N__29768;
    wire N__29767;
    wire N__29766;
    wire N__29765;
    wire N__29764;
    wire N__29761;
    wire N__29758;
    wire N__29753;
    wire N__29750;
    wire N__29747;
    wire N__29744;
    wire N__29741;
    wire N__29730;
    wire N__29727;
    wire N__29724;
    wire N__29721;
    wire N__29718;
    wire N__29717;
    wire N__29714;
    wire N__29711;
    wire N__29706;
    wire N__29703;
    wire N__29700;
    wire N__29697;
    wire N__29694;
    wire N__29691;
    wire N__29688;
    wire N__29685;
    wire N__29682;
    wire N__29679;
    wire N__29676;
    wire N__29673;
    wire N__29670;
    wire N__29667;
    wire N__29664;
    wire N__29663;
    wire N__29662;
    wire N__29661;
    wire N__29660;
    wire N__29659;
    wire N__29658;
    wire N__29653;
    wire N__29652;
    wire N__29649;
    wire N__29644;
    wire N__29643;
    wire N__29642;
    wire N__29637;
    wire N__29634;
    wire N__29633;
    wire N__29630;
    wire N__29629;
    wire N__29628;
    wire N__29625;
    wire N__29624;
    wire N__29623;
    wire N__29622;
    wire N__29621;
    wire N__29620;
    wire N__29619;
    wire N__29618;
    wire N__29615;
    wire N__29610;
    wire N__29605;
    wire N__29604;
    wire N__29603;
    wire N__29602;
    wire N__29601;
    wire N__29600;
    wire N__29599;
    wire N__29598;
    wire N__29591;
    wire N__29590;
    wire N__29589;
    wire N__29588;
    wire N__29587;
    wire N__29584;
    wire N__29581;
    wire N__29572;
    wire N__29569;
    wire N__29564;
    wire N__29561;
    wire N__29556;
    wire N__29545;
    wire N__29540;
    wire N__29537;
    wire N__29528;
    wire N__29521;
    wire N__29502;
    wire N__29501;
    wire N__29498;
    wire N__29497;
    wire N__29494;
    wire N__29491;
    wire N__29488;
    wire N__29481;
    wire N__29480;
    wire N__29479;
    wire N__29476;
    wire N__29471;
    wire N__29466;
    wire N__29463;
    wire N__29460;
    wire N__29457;
    wire N__29456;
    wire N__29453;
    wire N__29452;
    wire N__29451;
    wire N__29450;
    wire N__29449;
    wire N__29448;
    wire N__29445;
    wire N__29444;
    wire N__29443;
    wire N__29440;
    wire N__29431;
    wire N__29428;
    wire N__29427;
    wire N__29426;
    wire N__29425;
    wire N__29422;
    wire N__29419;
    wire N__29418;
    wire N__29417;
    wire N__29414;
    wire N__29413;
    wire N__29406;
    wire N__29401;
    wire N__29398;
    wire N__29393;
    wire N__29392;
    wire N__29389;
    wire N__29386;
    wire N__29383;
    wire N__29380;
    wire N__29375;
    wire N__29372;
    wire N__29369;
    wire N__29366;
    wire N__29363;
    wire N__29358;
    wire N__29355;
    wire N__29352;
    wire N__29349;
    wire N__29344;
    wire N__29339;
    wire N__29334;
    wire N__29325;
    wire N__29322;
    wire N__29319;
    wire N__29318;
    wire N__29315;
    wire N__29312;
    wire N__29309;
    wire N__29308;
    wire N__29305;
    wire N__29302;
    wire N__29299;
    wire N__29298;
    wire N__29291;
    wire N__29290;
    wire N__29287;
    wire N__29284;
    wire N__29281;
    wire N__29274;
    wire N__29271;
    wire N__29268;
    wire N__29265;
    wire N__29262;
    wire N__29261;
    wire N__29258;
    wire N__29257;
    wire N__29254;
    wire N__29249;
    wire N__29244;
    wire N__29243;
    wire N__29242;
    wire N__29239;
    wire N__29236;
    wire N__29233;
    wire N__29230;
    wire N__29223;
    wire N__29220;
    wire N__29217;
    wire N__29214;
    wire N__29211;
    wire N__29208;
    wire N__29205;
    wire N__29202;
    wire N__29199;
    wire N__29196;
    wire N__29193;
    wire N__29190;
    wire N__29187;
    wire N__29184;
    wire N__29181;
    wire N__29178;
    wire N__29175;
    wire N__29174;
    wire N__29171;
    wire N__29170;
    wire N__29167;
    wire N__29164;
    wire N__29161;
    wire N__29154;
    wire N__29153;
    wire N__29152;
    wire N__29149;
    wire N__29146;
    wire N__29143;
    wire N__29140;
    wire N__29133;
    wire N__29130;
    wire N__29127;
    wire N__29124;
    wire N__29121;
    wire N__29118;
    wire N__29115;
    wire N__29112;
    wire N__29109;
    wire N__29108;
    wire N__29107;
    wire N__29104;
    wire N__29101;
    wire N__29098;
    wire N__29095;
    wire N__29088;
    wire N__29087;
    wire N__29084;
    wire N__29083;
    wire N__29080;
    wire N__29077;
    wire N__29074;
    wire N__29067;
    wire N__29064;
    wire N__29061;
    wire N__29058;
    wire N__29055;
    wire N__29054;
    wire N__29053;
    wire N__29050;
    wire N__29045;
    wire N__29040;
    wire N__29039;
    wire N__29038;
    wire N__29035;
    wire N__29032;
    wire N__29029;
    wire N__29026;
    wire N__29019;
    wire N__29016;
    wire N__29013;
    wire N__29010;
    wire N__29007;
    wire N__29004;
    wire N__29003;
    wire N__29002;
    wire N__28999;
    wire N__28996;
    wire N__28993;
    wire N__28992;
    wire N__28991;
    wire N__28990;
    wire N__28989;
    wire N__28988;
    wire N__28987;
    wire N__28986;
    wire N__28985;
    wire N__28980;
    wire N__28977;
    wire N__28976;
    wire N__28973;
    wire N__28972;
    wire N__28967;
    wire N__28962;
    wire N__28959;
    wire N__28956;
    wire N__28953;
    wire N__28952;
    wire N__28947;
    wire N__28944;
    wire N__28943;
    wire N__28940;
    wire N__28937;
    wire N__28934;
    wire N__28925;
    wire N__28922;
    wire N__28919;
    wire N__28916;
    wire N__28913;
    wire N__28912;
    wire N__28909;
    wire N__28904;
    wire N__28899;
    wire N__28892;
    wire N__28889;
    wire N__28882;
    wire N__28875;
    wire N__28874;
    wire N__28873;
    wire N__28872;
    wire N__28871;
    wire N__28870;
    wire N__28867;
    wire N__28866;
    wire N__28863;
    wire N__28862;
    wire N__28861;
    wire N__28858;
    wire N__28855;
    wire N__28854;
    wire N__28851;
    wire N__28848;
    wire N__28847;
    wire N__28844;
    wire N__28839;
    wire N__28834;
    wire N__28833;
    wire N__28830;
    wire N__28827;
    wire N__28824;
    wire N__28823;
    wire N__28820;
    wire N__28819;
    wire N__28816;
    wire N__28813;
    wire N__28808;
    wire N__28805;
    wire N__28802;
    wire N__28801;
    wire N__28800;
    wire N__28797;
    wire N__28794;
    wire N__28791;
    wire N__28788;
    wire N__28785;
    wire N__28782;
    wire N__28779;
    wire N__28776;
    wire N__28769;
    wire N__28766;
    wire N__28763;
    wire N__28760;
    wire N__28753;
    wire N__28748;
    wire N__28737;
    wire N__28728;
    wire N__28727;
    wire N__28726;
    wire N__28725;
    wire N__28724;
    wire N__28723;
    wire N__28720;
    wire N__28719;
    wire N__28716;
    wire N__28715;
    wire N__28712;
    wire N__28711;
    wire N__28708;
    wire N__28705;
    wire N__28704;
    wire N__28703;
    wire N__28700;
    wire N__28699;
    wire N__28696;
    wire N__28693;
    wire N__28690;
    wire N__28687;
    wire N__28686;
    wire N__28685;
    wire N__28684;
    wire N__28681;
    wire N__28678;
    wire N__28677;
    wire N__28674;
    wire N__28671;
    wire N__28668;
    wire N__28665;
    wire N__28662;
    wire N__28659;
    wire N__28654;
    wire N__28649;
    wire N__28642;
    wire N__28639;
    wire N__28636;
    wire N__28633;
    wire N__28630;
    wire N__28623;
    wire N__28620;
    wire N__28617;
    wire N__28610;
    wire N__28603;
    wire N__28598;
    wire N__28591;
    wire N__28584;
    wire N__28581;
    wire N__28580;
    wire N__28579;
    wire N__28578;
    wire N__28577;
    wire N__28576;
    wire N__28573;
    wire N__28572;
    wire N__28569;
    wire N__28566;
    wire N__28565;
    wire N__28560;
    wire N__28559;
    wire N__28558;
    wire N__28557;
    wire N__28554;
    wire N__28551;
    wire N__28548;
    wire N__28545;
    wire N__28542;
    wire N__28541;
    wire N__28538;
    wire N__28535;
    wire N__28532;
    wire N__28529;
    wire N__28528;
    wire N__28527;
    wire N__28524;
    wire N__28523;
    wire N__28520;
    wire N__28515;
    wire N__28510;
    wire N__28507;
    wire N__28506;
    wire N__28503;
    wire N__28496;
    wire N__28491;
    wire N__28488;
    wire N__28485;
    wire N__28482;
    wire N__28479;
    wire N__28476;
    wire N__28473;
    wire N__28470;
    wire N__28463;
    wire N__28458;
    wire N__28453;
    wire N__28444;
    wire N__28437;
    wire N__28436;
    wire N__28435;
    wire N__28432;
    wire N__28429;
    wire N__28426;
    wire N__28423;
    wire N__28416;
    wire N__28415;
    wire N__28412;
    wire N__28411;
    wire N__28408;
    wire N__28405;
    wire N__28402;
    wire N__28399;
    wire N__28396;
    wire N__28389;
    wire N__28386;
    wire N__28383;
    wire N__28380;
    wire N__28377;
    wire N__28374;
    wire N__28371;
    wire N__28368;
    wire N__28367;
    wire N__28366;
    wire N__28363;
    wire N__28360;
    wire N__28355;
    wire N__28350;
    wire N__28349;
    wire N__28348;
    wire N__28345;
    wire N__28342;
    wire N__28339;
    wire N__28332;
    wire N__28329;
    wire N__28326;
    wire N__28323;
    wire N__28320;
    wire N__28317;
    wire N__28314;
    wire N__28311;
    wire N__28308;
    wire N__28305;
    wire N__28304;
    wire N__28301;
    wire N__28300;
    wire N__28297;
    wire N__28294;
    wire N__28291;
    wire N__28288;
    wire N__28283;
    wire N__28280;
    wire N__28277;
    wire N__28274;
    wire N__28269;
    wire N__28266;
    wire N__28265;
    wire N__28262;
    wire N__28259;
    wire N__28258;
    wire N__28255;
    wire N__28252;
    wire N__28249;
    wire N__28246;
    wire N__28241;
    wire N__28236;
    wire N__28233;
    wire N__28230;
    wire N__28227;
    wire N__28226;
    wire N__28223;
    wire N__28222;
    wire N__28219;
    wire N__28216;
    wire N__28213;
    wire N__28210;
    wire N__28207;
    wire N__28204;
    wire N__28201;
    wire N__28198;
    wire N__28191;
    wire N__28190;
    wire N__28189;
    wire N__28186;
    wire N__28183;
    wire N__28180;
    wire N__28177;
    wire N__28174;
    wire N__28171;
    wire N__28168;
    wire N__28161;
    wire N__28158;
    wire N__28155;
    wire N__28152;
    wire N__28149;
    wire N__28146;
    wire N__28143;
    wire N__28140;
    wire N__28139;
    wire N__28138;
    wire N__28137;
    wire N__28134;
    wire N__28133;
    wire N__28132;
    wire N__28129;
    wire N__28128;
    wire N__28127;
    wire N__28126;
    wire N__28123;
    wire N__28118;
    wire N__28115;
    wire N__28112;
    wire N__28109;
    wire N__28106;
    wire N__28103;
    wire N__28102;
    wire N__28101;
    wire N__28098;
    wire N__28095;
    wire N__28092;
    wire N__28089;
    wire N__28084;
    wire N__28081;
    wire N__28078;
    wire N__28075;
    wire N__28072;
    wire N__28067;
    wire N__28062;
    wire N__28059;
    wire N__28044;
    wire N__28043;
    wire N__28042;
    wire N__28039;
    wire N__28036;
    wire N__28033;
    wire N__28028;
    wire N__28025;
    wire N__28022;
    wire N__28017;
    wire N__28016;
    wire N__28015;
    wire N__28014;
    wire N__28013;
    wire N__28012;
    wire N__28009;
    wire N__28008;
    wire N__28005;
    wire N__28000;
    wire N__27997;
    wire N__27996;
    wire N__27993;
    wire N__27990;
    wire N__27989;
    wire N__27986;
    wire N__27983;
    wire N__27978;
    wire N__27977;
    wire N__27976;
    wire N__27973;
    wire N__27970;
    wire N__27967;
    wire N__27964;
    wire N__27961;
    wire N__27958;
    wire N__27955;
    wire N__27952;
    wire N__27949;
    wire N__27946;
    wire N__27941;
    wire N__27936;
    wire N__27931;
    wire N__27918;
    wire N__27917;
    wire N__27914;
    wire N__27913;
    wire N__27910;
    wire N__27907;
    wire N__27904;
    wire N__27901;
    wire N__27898;
    wire N__27895;
    wire N__27892;
    wire N__27889;
    wire N__27884;
    wire N__27879;
    wire N__27878;
    wire N__27875;
    wire N__27874;
    wire N__27871;
    wire N__27868;
    wire N__27865;
    wire N__27860;
    wire N__27857;
    wire N__27854;
    wire N__27851;
    wire N__27846;
    wire N__27843;
    wire N__27842;
    wire N__27841;
    wire N__27838;
    wire N__27835;
    wire N__27832;
    wire N__27829;
    wire N__27824;
    wire N__27819;
    wire N__27816;
    wire N__27813;
    wire N__27812;
    wire N__27809;
    wire N__27806;
    wire N__27803;
    wire N__27800;
    wire N__27797;
    wire N__27796;
    wire N__27793;
    wire N__27790;
    wire N__27787;
    wire N__27780;
    wire N__27777;
    wire N__27774;
    wire N__27771;
    wire N__27768;
    wire N__27765;
    wire N__27762;
    wire N__27759;
    wire N__27756;
    wire N__27753;
    wire N__27750;
    wire N__27747;
    wire N__27744;
    wire N__27741;
    wire N__27740;
    wire N__27737;
    wire N__27734;
    wire N__27731;
    wire N__27728;
    wire N__27725;
    wire N__27724;
    wire N__27721;
    wire N__27718;
    wire N__27715;
    wire N__27708;
    wire N__27705;
    wire N__27704;
    wire N__27701;
    wire N__27700;
    wire N__27697;
    wire N__27694;
    wire N__27691;
    wire N__27688;
    wire N__27685;
    wire N__27682;
    wire N__27679;
    wire N__27674;
    wire N__27669;
    wire N__27666;
    wire N__27663;
    wire N__27660;
    wire N__27657;
    wire N__27654;
    wire N__27651;
    wire N__27648;
    wire N__27645;
    wire N__27644;
    wire N__27641;
    wire N__27640;
    wire N__27637;
    wire N__27634;
    wire N__27631;
    wire N__27624;
    wire N__27621;
    wire N__27618;
    wire N__27615;
    wire N__27612;
    wire N__27609;
    wire N__27606;
    wire N__27603;
    wire N__27600;
    wire N__27599;
    wire N__27596;
    wire N__27595;
    wire N__27592;
    wire N__27589;
    wire N__27586;
    wire N__27583;
    wire N__27580;
    wire N__27577;
    wire N__27570;
    wire N__27569;
    wire N__27566;
    wire N__27565;
    wire N__27562;
    wire N__27559;
    wire N__27556;
    wire N__27553;
    wire N__27548;
    wire N__27543;
    wire N__27540;
    wire N__27537;
    wire N__27534;
    wire N__27531;
    wire N__27528;
    wire N__27527;
    wire N__27524;
    wire N__27521;
    wire N__27518;
    wire N__27517;
    wire N__27514;
    wire N__27511;
    wire N__27508;
    wire N__27501;
    wire N__27498;
    wire N__27495;
    wire N__27492;
    wire N__27489;
    wire N__27486;
    wire N__27483;
    wire N__27480;
    wire N__27477;
    wire N__27474;
    wire N__27473;
    wire N__27472;
    wire N__27469;
    wire N__27464;
    wire N__27459;
    wire N__27456;
    wire N__27453;
    wire N__27452;
    wire N__27451;
    wire N__27446;
    wire N__27445;
    wire N__27444;
    wire N__27443;
    wire N__27442;
    wire N__27441;
    wire N__27440;
    wire N__27439;
    wire N__27436;
    wire N__27433;
    wire N__27432;
    wire N__27431;
    wire N__27428;
    wire N__27427;
    wire N__27424;
    wire N__27423;
    wire N__27422;
    wire N__27419;
    wire N__27416;
    wire N__27415;
    wire N__27412;
    wire N__27409;
    wire N__27404;
    wire N__27401;
    wire N__27398;
    wire N__27393;
    wire N__27386;
    wire N__27377;
    wire N__27372;
    wire N__27369;
    wire N__27354;
    wire N__27353;
    wire N__27352;
    wire N__27351;
    wire N__27348;
    wire N__27347;
    wire N__27346;
    wire N__27345;
    wire N__27344;
    wire N__27343;
    wire N__27342;
    wire N__27339;
    wire N__27338;
    wire N__27333;
    wire N__27332;
    wire N__27331;
    wire N__27330;
    wire N__27327;
    wire N__27320;
    wire N__27313;
    wire N__27308;
    wire N__27305;
    wire N__27298;
    wire N__27285;
    wire N__27282;
    wire N__27279;
    wire N__27276;
    wire N__27273;
    wire N__27270;
    wire N__27267;
    wire N__27264;
    wire N__27263;
    wire N__27260;
    wire N__27259;
    wire N__27256;
    wire N__27253;
    wire N__27250;
    wire N__27247;
    wire N__27244;
    wire N__27241;
    wire N__27234;
    wire N__27231;
    wire N__27228;
    wire N__27225;
    wire N__27222;
    wire N__27221;
    wire N__27220;
    wire N__27217;
    wire N__27214;
    wire N__27211;
    wire N__27206;
    wire N__27203;
    wire N__27200;
    wire N__27195;
    wire N__27192;
    wire N__27189;
    wire N__27186;
    wire N__27183;
    wire N__27180;
    wire N__27179;
    wire N__27178;
    wire N__27175;
    wire N__27172;
    wire N__27169;
    wire N__27166;
    wire N__27159;
    wire N__27156;
    wire N__27153;
    wire N__27150;
    wire N__27147;
    wire N__27144;
    wire N__27141;
    wire N__27138;
    wire N__27135;
    wire N__27134;
    wire N__27131;
    wire N__27128;
    wire N__27125;
    wire N__27120;
    wire N__27117;
    wire N__27114;
    wire N__27111;
    wire N__27108;
    wire N__27105;
    wire N__27102;
    wire N__27099;
    wire N__27096;
    wire N__27093;
    wire N__27090;
    wire N__27087;
    wire N__27084;
    wire N__27081;
    wire N__27078;
    wire N__27075;
    wire N__27072;
    wire N__27069;
    wire N__27066;
    wire N__27063;
    wire N__27060;
    wire N__27057;
    wire N__27054;
    wire N__27053;
    wire N__27052;
    wire N__27049;
    wire N__27046;
    wire N__27043;
    wire N__27036;
    wire N__27033;
    wire N__27030;
    wire N__27027;
    wire N__27024;
    wire N__27021;
    wire N__27018;
    wire N__27015;
    wire N__27012;
    wire N__27009;
    wire N__27008;
    wire N__27007;
    wire N__27004;
    wire N__26999;
    wire N__26994;
    wire N__26993;
    wire N__26992;
    wire N__26989;
    wire N__26986;
    wire N__26983;
    wire N__26976;
    wire N__26975;
    wire N__26974;
    wire N__26967;
    wire N__26964;
    wire N__26961;
    wire N__26958;
    wire N__26955;
    wire N__26954;
    wire N__26953;
    wire N__26952;
    wire N__26949;
    wire N__26946;
    wire N__26943;
    wire N__26940;
    wire N__26935;
    wire N__26934;
    wire N__26931;
    wire N__26928;
    wire N__26925;
    wire N__26922;
    wire N__26919;
    wire N__26916;
    wire N__26911;
    wire N__26904;
    wire N__26903;
    wire N__26898;
    wire N__26895;
    wire N__26892;
    wire N__26889;
    wire N__26888;
    wire N__26887;
    wire N__26884;
    wire N__26883;
    wire N__26874;
    wire N__26871;
    wire N__26870;
    wire N__26869;
    wire N__26868;
    wire N__26859;
    wire N__26856;
    wire N__26855;
    wire N__26852;
    wire N__26849;
    wire N__26846;
    wire N__26841;
    wire N__26838;
    wire N__26835;
    wire N__26834;
    wire N__26833;
    wire N__26830;
    wire N__26827;
    wire N__26824;
    wire N__26821;
    wire N__26814;
    wire N__26813;
    wire N__26812;
    wire N__26809;
    wire N__26806;
    wire N__26803;
    wire N__26800;
    wire N__26793;
    wire N__26790;
    wire N__26787;
    wire N__26784;
    wire N__26781;
    wire N__26778;
    wire N__26775;
    wire N__26772;
    wire N__26769;
    wire N__26766;
    wire N__26763;
    wire N__26760;
    wire N__26757;
    wire N__26754;
    wire N__26751;
    wire N__26750;
    wire N__26749;
    wire N__26748;
    wire N__26747;
    wire N__26746;
    wire N__26743;
    wire N__26740;
    wire N__26737;
    wire N__26732;
    wire N__26729;
    wire N__26726;
    wire N__26715;
    wire N__26712;
    wire N__26709;
    wire N__26706;
    wire N__26705;
    wire N__26704;
    wire N__26699;
    wire N__26696;
    wire N__26693;
    wire N__26688;
    wire N__26685;
    wire N__26684;
    wire N__26683;
    wire N__26680;
    wire N__26677;
    wire N__26674;
    wire N__26669;
    wire N__26664;
    wire N__26663;
    wire N__26662;
    wire N__26659;
    wire N__26654;
    wire N__26649;
    wire N__26646;
    wire N__26643;
    wire N__26640;
    wire N__26637;
    wire N__26634;
    wire N__26631;
    wire N__26628;
    wire N__26625;
    wire N__26622;
    wire N__26619;
    wire N__26618;
    wire N__26617;
    wire N__26614;
    wire N__26609;
    wire N__26604;
    wire N__26601;
    wire N__26598;
    wire N__26595;
    wire N__26592;
    wire N__26589;
    wire N__26586;
    wire N__26583;
    wire N__26580;
    wire N__26577;
    wire N__26574;
    wire N__26571;
    wire N__26568;
    wire N__26567;
    wire N__26564;
    wire N__26563;
    wire N__26560;
    wire N__26555;
    wire N__26550;
    wire N__26549;
    wire N__26548;
    wire N__26545;
    wire N__26542;
    wire N__26539;
    wire N__26536;
    wire N__26533;
    wire N__26526;
    wire N__26523;
    wire N__26520;
    wire N__26517;
    wire N__26514;
    wire N__26511;
    wire N__26508;
    wire N__26505;
    wire N__26502;
    wire N__26499;
    wire N__26496;
    wire N__26493;
    wire N__26492;
    wire N__26491;
    wire N__26486;
    wire N__26483;
    wire N__26480;
    wire N__26475;
    wire N__26472;
    wire N__26469;
    wire N__26466;
    wire N__26463;
    wire N__26460;
    wire N__26457;
    wire N__26454;
    wire N__26451;
    wire N__26448;
    wire N__26445;
    wire N__26442;
    wire N__26439;
    wire N__26436;
    wire N__26433;
    wire N__26432;
    wire N__26429;
    wire N__26428;
    wire N__26425;
    wire N__26422;
    wire N__26419;
    wire N__26412;
    wire N__26409;
    wire N__26406;
    wire N__26403;
    wire N__26402;
    wire N__26401;
    wire N__26398;
    wire N__26393;
    wire N__26388;
    wire N__26385;
    wire N__26382;
    wire N__26379;
    wire N__26376;
    wire N__26375;
    wire N__26374;
    wire N__26371;
    wire N__26368;
    wire N__26365;
    wire N__26362;
    wire N__26359;
    wire N__26356;
    wire N__26353;
    wire N__26350;
    wire N__26345;
    wire N__26340;
    wire N__26337;
    wire N__26336;
    wire N__26333;
    wire N__26330;
    wire N__26329;
    wire N__26326;
    wire N__26323;
    wire N__26320;
    wire N__26317;
    wire N__26312;
    wire N__26309;
    wire N__26304;
    wire N__26303;
    wire N__26300;
    wire N__26297;
    wire N__26294;
    wire N__26291;
    wire N__26288;
    wire N__26287;
    wire N__26284;
    wire N__26281;
    wire N__26278;
    wire N__26271;
    wire N__26270;
    wire N__26267;
    wire N__26264;
    wire N__26261;
    wire N__26258;
    wire N__26257;
    wire N__26252;
    wire N__26249;
    wire N__26244;
    wire N__26241;
    wire N__26238;
    wire N__26235;
    wire N__26232;
    wire N__26229;
    wire N__26226;
    wire N__26223;
    wire N__26220;
    wire N__26217;
    wire N__26214;
    wire N__26211;
    wire N__26208;
    wire N__26205;
    wire N__26202;
    wire N__26199;
    wire N__26196;
    wire N__26193;
    wire N__26190;
    wire N__26187;
    wire N__26184;
    wire N__26183;
    wire N__26182;
    wire N__26181;
    wire N__26180;
    wire N__26179;
    wire N__26178;
    wire N__26163;
    wire N__26160;
    wire N__26157;
    wire N__26156;
    wire N__26155;
    wire N__26154;
    wire N__26153;
    wire N__26152;
    wire N__26151;
    wire N__26136;
    wire N__26133;
    wire N__26130;
    wire N__26127;
    wire N__26124;
    wire N__26121;
    wire N__26118;
    wire N__26115;
    wire N__26112;
    wire N__26109;
    wire N__26108;
    wire N__26107;
    wire N__26104;
    wire N__26101;
    wire N__26098;
    wire N__26093;
    wire N__26090;
    wire N__26087;
    wire N__26084;
    wire N__26079;
    wire N__26076;
    wire N__26073;
    wire N__26070;
    wire N__26067;
    wire N__26064;
    wire N__26061;
    wire N__26058;
    wire N__26055;
    wire N__26054;
    wire N__26053;
    wire N__26052;
    wire N__26047;
    wire N__26044;
    wire N__26043;
    wire N__26042;
    wire N__26041;
    wire N__26040;
    wire N__26039;
    wire N__26038;
    wire N__26037;
    wire N__26034;
    wire N__26031;
    wire N__26028;
    wire N__26025;
    wire N__26022;
    wire N__26015;
    wire N__26014;
    wire N__26013;
    wire N__26012;
    wire N__26011;
    wire N__26008;
    wire N__26005;
    wire N__26004;
    wire N__26001;
    wire N__25994;
    wire N__25991;
    wire N__25988;
    wire N__25983;
    wire N__25980;
    wire N__25977;
    wire N__25976;
    wire N__25975;
    wire N__25974;
    wire N__25973;
    wire N__25972;
    wire N__25971;
    wire N__25970;
    wire N__25969;
    wire N__25966;
    wire N__25961;
    wire N__25956;
    wire N__25951;
    wire N__25946;
    wire N__25943;
    wire N__25936;
    wire N__25935;
    wire N__25932;
    wire N__25929;
    wire N__25928;
    wire N__25927;
    wire N__25924;
    wire N__25921;
    wire N__25920;
    wire N__25919;
    wire N__25918;
    wire N__25917;
    wire N__25914;
    wire N__25907;
    wire N__25902;
    wire N__25897;
    wire N__25888;
    wire N__25877;
    wire N__25872;
    wire N__25857;
    wire N__25854;
    wire N__25851;
    wire N__25848;
    wire N__25845;
    wire N__25842;
    wire N__25841;
    wire N__25838;
    wire N__25835;
    wire N__25834;
    wire N__25831;
    wire N__25828;
    wire N__25825;
    wire N__25822;
    wire N__25819;
    wire N__25816;
    wire N__25813;
    wire N__25806;
    wire N__25803;
    wire N__25802;
    wire N__25801;
    wire N__25800;
    wire N__25799;
    wire N__25798;
    wire N__25797;
    wire N__25796;
    wire N__25795;
    wire N__25792;
    wire N__25789;
    wire N__25786;
    wire N__25779;
    wire N__25778;
    wire N__25773;
    wire N__25772;
    wire N__25769;
    wire N__25764;
    wire N__25761;
    wire N__25758;
    wire N__25757;
    wire N__25756;
    wire N__25753;
    wire N__25750;
    wire N__25747;
    wire N__25744;
    wire N__25739;
    wire N__25736;
    wire N__25735;
    wire N__25734;
    wire N__25733;
    wire N__25732;
    wire N__25731;
    wire N__25730;
    wire N__25729;
    wire N__25728;
    wire N__25727;
    wire N__25726;
    wire N__25725;
    wire N__25724;
    wire N__25723;
    wire N__25722;
    wire N__25721;
    wire N__25720;
    wire N__25717;
    wire N__25716;
    wire N__25715;
    wire N__25712;
    wire N__25707;
    wire N__25702;
    wire N__25697;
    wire N__25680;
    wire N__25669;
    wire N__25656;
    wire N__25641;
    wire N__25638;
    wire N__25635;
    wire N__25632;
    wire N__25629;
    wire N__25626;
    wire N__25623;
    wire N__25620;
    wire N__25617;
    wire N__25614;
    wire N__25611;
    wire N__25608;
    wire N__25607;
    wire N__25604;
    wire N__25601;
    wire N__25598;
    wire N__25597;
    wire N__25594;
    wire N__25591;
    wire N__25588;
    wire N__25583;
    wire N__25580;
    wire N__25575;
    wire N__25572;
    wire N__25569;
    wire N__25568;
    wire N__25567;
    wire N__25564;
    wire N__25561;
    wire N__25558;
    wire N__25555;
    wire N__25550;
    wire N__25545;
    wire N__25544;
    wire N__25541;
    wire N__25538;
    wire N__25535;
    wire N__25532;
    wire N__25531;
    wire N__25526;
    wire N__25523;
    wire N__25518;
    wire N__25515;
    wire N__25514;
    wire N__25511;
    wire N__25508;
    wire N__25507;
    wire N__25504;
    wire N__25501;
    wire N__25498;
    wire N__25495;
    wire N__25490;
    wire N__25485;
    wire N__25482;
    wire N__25481;
    wire N__25480;
    wire N__25477;
    wire N__25474;
    wire N__25471;
    wire N__25468;
    wire N__25463;
    wire N__25460;
    wire N__25455;
    wire N__25452;
    wire N__25449;
    wire N__25446;
    wire N__25443;
    wire N__25442;
    wire N__25439;
    wire N__25438;
    wire N__25435;
    wire N__25432;
    wire N__25429;
    wire N__25424;
    wire N__25419;
    wire N__25418;
    wire N__25415;
    wire N__25414;
    wire N__25411;
    wire N__25408;
    wire N__25405;
    wire N__25400;
    wire N__25397;
    wire N__25392;
    wire N__25391;
    wire N__25388;
    wire N__25387;
    wire N__25384;
    wire N__25381;
    wire N__25378;
    wire N__25375;
    wire N__25370;
    wire N__25367;
    wire N__25364;
    wire N__25359;
    wire N__25356;
    wire N__25353;
    wire N__25350;
    wire N__25349;
    wire N__25348;
    wire N__25345;
    wire N__25342;
    wire N__25339;
    wire N__25336;
    wire N__25331;
    wire N__25328;
    wire N__25323;
    wire N__25320;
    wire N__25317;
    wire N__25314;
    wire N__25311;
    wire N__25310;
    wire N__25307;
    wire N__25304;
    wire N__25303;
    wire N__25300;
    wire N__25297;
    wire N__25294;
    wire N__25291;
    wire N__25286;
    wire N__25281;
    wire N__25280;
    wire N__25277;
    wire N__25274;
    wire N__25271;
    wire N__25268;
    wire N__25267;
    wire N__25262;
    wire N__25259;
    wire N__25254;
    wire N__25251;
    wire N__25248;
    wire N__25245;
    wire N__25242;
    wire N__25239;
    wire N__25236;
    wire N__25233;
    wire N__25230;
    wire N__25227;
    wire N__25224;
    wire N__25221;
    wire N__25218;
    wire N__25215;
    wire N__25214;
    wire N__25211;
    wire N__25208;
    wire N__25205;
    wire N__25202;
    wire N__25197;
    wire N__25194;
    wire N__25191;
    wire N__25188;
    wire N__25185;
    wire N__25182;
    wire N__25179;
    wire N__25176;
    wire N__25173;
    wire N__25170;
    wire N__25167;
    wire N__25164;
    wire N__25161;
    wire N__25158;
    wire N__25155;
    wire N__25152;
    wire N__25149;
    wire N__25146;
    wire N__25143;
    wire N__25140;
    wire N__25137;
    wire N__25134;
    wire N__25131;
    wire N__25128;
    wire N__25125;
    wire N__25122;
    wire N__25119;
    wire N__25116;
    wire N__25115;
    wire N__25112;
    wire N__25109;
    wire N__25108;
    wire N__25105;
    wire N__25102;
    wire N__25099;
    wire N__25096;
    wire N__25089;
    wire N__25088;
    wire N__25087;
    wire N__25084;
    wire N__25081;
    wire N__25078;
    wire N__25075;
    wire N__25072;
    wire N__25069;
    wire N__25062;
    wire N__25059;
    wire N__25056;
    wire N__25053;
    wire N__25050;
    wire N__25047;
    wire N__25044;
    wire N__25041;
    wire N__25038;
    wire N__25035;
    wire N__25032;
    wire N__25029;
    wire N__25026;
    wire N__25023;
    wire N__25020;
    wire N__25017;
    wire N__25014;
    wire N__25011;
    wire N__25008;
    wire N__25005;
    wire N__25002;
    wire N__24999;
    wire N__24996;
    wire N__24993;
    wire N__24990;
    wire N__24987;
    wire N__24984;
    wire N__24981;
    wire N__24978;
    wire N__24975;
    wire N__24972;
    wire N__24969;
    wire N__24966;
    wire N__24963;
    wire N__24962;
    wire N__24959;
    wire N__24956;
    wire N__24951;
    wire N__24948;
    wire N__24945;
    wire N__24942;
    wire N__24939;
    wire N__24936;
    wire N__24933;
    wire N__24930;
    wire N__24927;
    wire N__24924;
    wire N__24921;
    wire N__24918;
    wire N__24915;
    wire N__24914;
    wire N__24911;
    wire N__24910;
    wire N__24907;
    wire N__24904;
    wire N__24901;
    wire N__24894;
    wire N__24891;
    wire N__24888;
    wire N__24885;
    wire N__24882;
    wire N__24879;
    wire N__24876;
    wire N__24873;
    wire N__24870;
    wire N__24867;
    wire N__24864;
    wire N__24861;
    wire N__24858;
    wire N__24855;
    wire N__24852;
    wire N__24849;
    wire N__24846;
    wire N__24843;
    wire N__24840;
    wire N__24837;
    wire N__24834;
    wire N__24833;
    wire N__24832;
    wire N__24829;
    wire N__24826;
    wire N__24823;
    wire N__24820;
    wire N__24813;
    wire N__24810;
    wire N__24807;
    wire N__24804;
    wire N__24801;
    wire N__24798;
    wire N__24797;
    wire N__24796;
    wire N__24793;
    wire N__24788;
    wire N__24783;
    wire N__24780;
    wire N__24777;
    wire N__24776;
    wire N__24775;
    wire N__24772;
    wire N__24769;
    wire N__24766;
    wire N__24763;
    wire N__24760;
    wire N__24753;
    wire N__24750;
    wire N__24749;
    wire N__24746;
    wire N__24745;
    wire N__24742;
    wire N__24739;
    wire N__24736;
    wire N__24729;
    wire N__24726;
    wire N__24723;
    wire N__24720;
    wire N__24717;
    wire N__24714;
    wire N__24711;
    wire N__24708;
    wire N__24705;
    wire N__24702;
    wire N__24699;
    wire N__24696;
    wire N__24695;
    wire N__24694;
    wire N__24691;
    wire N__24688;
    wire N__24685;
    wire N__24678;
    wire N__24675;
    wire N__24674;
    wire N__24673;
    wire N__24670;
    wire N__24667;
    wire N__24662;
    wire N__24657;
    wire N__24654;
    wire N__24653;
    wire N__24652;
    wire N__24649;
    wire N__24644;
    wire N__24639;
    wire N__24636;
    wire N__24635;
    wire N__24634;
    wire N__24629;
    wire N__24626;
    wire N__24621;
    wire N__24620;
    wire N__24615;
    wire N__24612;
    wire N__24611;
    wire N__24608;
    wire N__24605;
    wire N__24604;
    wire N__24603;
    wire N__24594;
    wire N__24591;
    wire N__24590;
    wire N__24589;
    wire N__24588;
    wire N__24579;
    wire N__24576;
    wire N__24573;
    wire N__24570;
    wire N__24567;
    wire N__24564;
    wire N__24561;
    wire N__24558;
    wire N__24557;
    wire N__24556;
    wire N__24553;
    wire N__24552;
    wire N__24549;
    wire N__24546;
    wire N__24543;
    wire N__24540;
    wire N__24539;
    wire N__24536;
    wire N__24533;
    wire N__24530;
    wire N__24527;
    wire N__24524;
    wire N__24521;
    wire N__24518;
    wire N__24513;
    wire N__24510;
    wire N__24507;
    wire N__24498;
    wire N__24495;
    wire N__24492;
    wire N__24489;
    wire N__24486;
    wire N__24485;
    wire N__24482;
    wire N__24479;
    wire N__24474;
    wire N__24473;
    wire N__24470;
    wire N__24467;
    wire N__24462;
    wire N__24461;
    wire N__24458;
    wire N__24455;
    wire N__24450;
    wire N__24449;
    wire N__24446;
    wire N__24443;
    wire N__24438;
    wire N__24437;
    wire N__24434;
    wire N__24431;
    wire N__24426;
    wire N__24425;
    wire N__24422;
    wire N__24419;
    wire N__24414;
    wire N__24411;
    wire N__24410;
    wire N__24407;
    wire N__24406;
    wire N__24403;
    wire N__24400;
    wire N__24397;
    wire N__24394;
    wire N__24389;
    wire N__24386;
    wire N__24383;
    wire N__24380;
    wire N__24375;
    wire N__24374;
    wire N__24371;
    wire N__24368;
    wire N__24367;
    wire N__24364;
    wire N__24361;
    wire N__24358;
    wire N__24355;
    wire N__24352;
    wire N__24349;
    wire N__24346;
    wire N__24341;
    wire N__24336;
    wire N__24335;
    wire N__24332;
    wire N__24329;
    wire N__24326;
    wire N__24323;
    wire N__24320;
    wire N__24315;
    wire N__24314;
    wire N__24311;
    wire N__24308;
    wire N__24305;
    wire N__24302;
    wire N__24299;
    wire N__24294;
    wire N__24291;
    wire N__24290;
    wire N__24287;
    wire N__24284;
    wire N__24281;
    wire N__24276;
    wire N__24273;
    wire N__24270;
    wire N__24269;
    wire N__24266;
    wire N__24263;
    wire N__24260;
    wire N__24257;
    wire N__24252;
    wire N__24249;
    wire N__24246;
    wire N__24243;
    wire N__24242;
    wire N__24239;
    wire N__24236;
    wire N__24233;
    wire N__24228;
    wire N__24227;
    wire N__24224;
    wire N__24221;
    wire N__24218;
    wire N__24213;
    wire N__24210;
    wire N__24209;
    wire N__24208;
    wire N__24205;
    wire N__24202;
    wire N__24201;
    wire N__24200;
    wire N__24199;
    wire N__24198;
    wire N__24197;
    wire N__24196;
    wire N__24183;
    wire N__24182;
    wire N__24181;
    wire N__24180;
    wire N__24179;
    wire N__24178;
    wire N__24175;
    wire N__24174;
    wire N__24173;
    wire N__24170;
    wire N__24167;
    wire N__24164;
    wire N__24157;
    wire N__24144;
    wire N__24135;
    wire N__24132;
    wire N__24129;
    wire N__24128;
    wire N__24125;
    wire N__24122;
    wire N__24121;
    wire N__24118;
    wire N__24115;
    wire N__24112;
    wire N__24109;
    wire N__24102;
    wire N__24101;
    wire N__24100;
    wire N__24099;
    wire N__24098;
    wire N__24097;
    wire N__24096;
    wire N__24095;
    wire N__24092;
    wire N__24087;
    wire N__24086;
    wire N__24085;
    wire N__24084;
    wire N__24081;
    wire N__24080;
    wire N__24077;
    wire N__24072;
    wire N__24069;
    wire N__24066;
    wire N__24063;
    wire N__24060;
    wire N__24059;
    wire N__24056;
    wire N__24053;
    wire N__24052;
    wire N__24051;
    wire N__24050;
    wire N__24045;
    wire N__24042;
    wire N__24037;
    wire N__24032;
    wire N__24029;
    wire N__24028;
    wire N__24027;
    wire N__24026;
    wire N__24025;
    wire N__24024;
    wire N__24023;
    wire N__24022;
    wire N__24021;
    wire N__24018;
    wire N__24011;
    wire N__24010;
    wire N__24009;
    wire N__24008;
    wire N__24007;
    wire N__24006;
    wire N__24005;
    wire N__24004;
    wire N__24001;
    wire N__23998;
    wire N__23993;
    wire N__23990;
    wire N__23985;
    wire N__23968;
    wire N__23963;
    wire N__23950;
    wire N__23947;
    wire N__23928;
    wire N__23925;
    wire N__23922;
    wire N__23919;
    wire N__23918;
    wire N__23917;
    wire N__23914;
    wire N__23911;
    wire N__23908;
    wire N__23905;
    wire N__23898;
    wire N__23897;
    wire N__23894;
    wire N__23891;
    wire N__23890;
    wire N__23887;
    wire N__23884;
    wire N__23881;
    wire N__23878;
    wire N__23873;
    wire N__23868;
    wire N__23865;
    wire N__23862;
    wire N__23859;
    wire N__23858;
    wire N__23855;
    wire N__23854;
    wire N__23851;
    wire N__23848;
    wire N__23845;
    wire N__23838;
    wire N__23835;
    wire N__23834;
    wire N__23831;
    wire N__23828;
    wire N__23827;
    wire N__23822;
    wire N__23819;
    wire N__23816;
    wire N__23811;
    wire N__23808;
    wire N__23807;
    wire N__23804;
    wire N__23801;
    wire N__23800;
    wire N__23795;
    wire N__23792;
    wire N__23787;
    wire N__23784;
    wire N__23783;
    wire N__23782;
    wire N__23779;
    wire N__23776;
    wire N__23773;
    wire N__23770;
    wire N__23767;
    wire N__23760;
    wire N__23757;
    wire N__23754;
    wire N__23751;
    wire N__23748;
    wire N__23745;
    wire N__23742;
    wire N__23741;
    wire N__23738;
    wire N__23735;
    wire N__23734;
    wire N__23729;
    wire N__23726;
    wire N__23721;
    wire N__23718;
    wire N__23717;
    wire N__23714;
    wire N__23711;
    wire N__23710;
    wire N__23707;
    wire N__23704;
    wire N__23701;
    wire N__23696;
    wire N__23693;
    wire N__23688;
    wire N__23685;
    wire N__23682;
    wire N__23679;
    wire N__23676;
    wire N__23673;
    wire N__23670;
    wire N__23667;
    wire N__23664;
    wire N__23661;
    wire N__23658;
    wire N__23655;
    wire N__23652;
    wire N__23649;
    wire N__23646;
    wire N__23643;
    wire N__23640;
    wire N__23637;
    wire N__23634;
    wire N__23631;
    wire N__23628;
    wire N__23625;
    wire N__23624;
    wire N__23623;
    wire N__23622;
    wire N__23619;
    wire N__23618;
    wire N__23615;
    wire N__23614;
    wire N__23613;
    wire N__23612;
    wire N__23611;
    wire N__23610;
    wire N__23599;
    wire N__23596;
    wire N__23595;
    wire N__23592;
    wire N__23589;
    wire N__23588;
    wire N__23585;
    wire N__23582;
    wire N__23581;
    wire N__23580;
    wire N__23579;
    wire N__23576;
    wire N__23563;
    wire N__23554;
    wire N__23547;
    wire N__23544;
    wire N__23541;
    wire N__23538;
    wire N__23535;
    wire N__23532;
    wire N__23529;
    wire N__23526;
    wire N__23523;
    wire N__23520;
    wire N__23517;
    wire N__23514;
    wire N__23511;
    wire N__23508;
    wire N__23505;
    wire N__23502;
    wire N__23501;
    wire N__23496;
    wire N__23493;
    wire N__23492;
    wire N__23491;
    wire N__23484;
    wire N__23481;
    wire N__23478;
    wire N__23475;
    wire N__23472;
    wire N__23469;
    wire N__23466;
    wire N__23463;
    wire N__23460;
    wire N__23459;
    wire N__23458;
    wire N__23455;
    wire N__23452;
    wire N__23451;
    wire N__23450;
    wire N__23449;
    wire N__23448;
    wire N__23445;
    wire N__23444;
    wire N__23441;
    wire N__23438;
    wire N__23435;
    wire N__23430;
    wire N__23429;
    wire N__23428;
    wire N__23425;
    wire N__23422;
    wire N__23419;
    wire N__23410;
    wire N__23405;
    wire N__23402;
    wire N__23397;
    wire N__23392;
    wire N__23391;
    wire N__23388;
    wire N__23385;
    wire N__23382;
    wire N__23379;
    wire N__23370;
    wire N__23367;
    wire N__23366;
    wire N__23363;
    wire N__23362;
    wire N__23359;
    wire N__23356;
    wire N__23353;
    wire N__23350;
    wire N__23345;
    wire N__23340;
    wire N__23337;
    wire N__23334;
    wire N__23331;
    wire N__23328;
    wire N__23325;
    wire N__23322;
    wire N__23319;
    wire N__23316;
    wire N__23313;
    wire N__23310;
    wire N__23307;
    wire N__23304;
    wire N__23301;
    wire N__23298;
    wire N__23295;
    wire N__23292;
    wire N__23289;
    wire N__23286;
    wire N__23283;
    wire N__23280;
    wire N__23277;
    wire N__23274;
    wire N__23271;
    wire N__23268;
    wire N__23265;
    wire N__23264;
    wire N__23263;
    wire N__23260;
    wire N__23257;
    wire N__23254;
    wire N__23251;
    wire N__23246;
    wire N__23241;
    wire N__23238;
    wire N__23235;
    wire N__23232;
    wire N__23231;
    wire N__23228;
    wire N__23225;
    wire N__23222;
    wire N__23217;
    wire N__23214;
    wire N__23211;
    wire N__23208;
    wire N__23205;
    wire N__23202;
    wire N__23199;
    wire N__23196;
    wire N__23195;
    wire N__23192;
    wire N__23189;
    wire N__23188;
    wire N__23183;
    wire N__23180;
    wire N__23175;
    wire N__23174;
    wire N__23171;
    wire N__23168;
    wire N__23167;
    wire N__23162;
    wire N__23159;
    wire N__23154;
    wire N__23151;
    wire N__23148;
    wire N__23145;
    wire N__23142;
    wire N__23139;
    wire N__23136;
    wire N__23133;
    wire N__23130;
    wire N__23129;
    wire N__23128;
    wire N__23125;
    wire N__23122;
    wire N__23119;
    wire N__23116;
    wire N__23109;
    wire N__23106;
    wire N__23103;
    wire N__23102;
    wire N__23099;
    wire N__23098;
    wire N__23095;
    wire N__23092;
    wire N__23089;
    wire N__23086;
    wire N__23083;
    wire N__23076;
    wire N__23073;
    wire N__23070;
    wire N__23067;
    wire N__23064;
    wire N__23061;
    wire N__23058;
    wire N__23055;
    wire N__23054;
    wire N__23053;
    wire N__23050;
    wire N__23047;
    wire N__23044;
    wire N__23041;
    wire N__23034;
    wire N__23031;
    wire N__23030;
    wire N__23027;
    wire N__23026;
    wire N__23023;
    wire N__23020;
    wire N__23017;
    wire N__23010;
    wire N__23007;
    wire N__23004;
    wire N__23001;
    wire N__22998;
    wire N__22995;
    wire N__22994;
    wire N__22993;
    wire N__22990;
    wire N__22985;
    wire N__22980;
    wire N__22979;
    wire N__22978;
    wire N__22975;
    wire N__22972;
    wire N__22965;
    wire N__22962;
    wire N__22959;
    wire N__22956;
    wire N__22953;
    wire N__22950;
    wire N__22947;
    wire N__22944;
    wire N__22941;
    wire N__22938;
    wire N__22935;
    wire N__22932;
    wire N__22929;
    wire N__22926;
    wire N__22923;
    wire N__22922;
    wire N__22919;
    wire N__22916;
    wire N__22911;
    wire N__22910;
    wire N__22907;
    wire N__22904;
    wire N__22899;
    wire N__22898;
    wire N__22895;
    wire N__22892;
    wire N__22887;
    wire N__22886;
    wire N__22883;
    wire N__22880;
    wire N__22875;
    wire N__22874;
    wire N__22871;
    wire N__22868;
    wire N__22863;
    wire N__22862;
    wire N__22861;
    wire N__22858;
    wire N__22855;
    wire N__22852;
    wire N__22845;
    wire N__22842;
    wire N__22839;
    wire N__22838;
    wire N__22835;
    wire N__22832;
    wire N__22829;
    wire N__22826;
    wire N__22823;
    wire N__22822;
    wire N__22819;
    wire N__22816;
    wire N__22813;
    wire N__22806;
    wire N__22805;
    wire N__22802;
    wire N__22799;
    wire N__22798;
    wire N__22797;
    wire N__22796;
    wire N__22795;
    wire N__22794;
    wire N__22793;
    wire N__22792;
    wire N__22791;
    wire N__22790;
    wire N__22789;
    wire N__22788;
    wire N__22787;
    wire N__22784;
    wire N__22783;
    wire N__22780;
    wire N__22777;
    wire N__22772;
    wire N__22765;
    wire N__22762;
    wire N__22759;
    wire N__22758;
    wire N__22757;
    wire N__22756;
    wire N__22755;
    wire N__22754;
    wire N__22753;
    wire N__22750;
    wire N__22743;
    wire N__22740;
    wire N__22737;
    wire N__22730;
    wire N__22723;
    wire N__22722;
    wire N__22721;
    wire N__22720;
    wire N__22719;
    wire N__22718;
    wire N__22717;
    wire N__22714;
    wire N__22711;
    wire N__22710;
    wire N__22707;
    wire N__22706;
    wire N__22705;
    wire N__22704;
    wire N__22701;
    wire N__22698;
    wire N__22695;
    wire N__22688;
    wire N__22681;
    wire N__22676;
    wire N__22667;
    wire N__22652;
    wire N__22635;
    wire N__22634;
    wire N__22633;
    wire N__22632;
    wire N__22631;
    wire N__22630;
    wire N__22627;
    wire N__22624;
    wire N__22621;
    wire N__22618;
    wire N__22615;
    wire N__22614;
    wire N__22611;
    wire N__22610;
    wire N__22609;
    wire N__22608;
    wire N__22607;
    wire N__22606;
    wire N__22605;
    wire N__22604;
    wire N__22599;
    wire N__22594;
    wire N__22587;
    wire N__22572;
    wire N__22563;
    wire N__22562;
    wire N__22559;
    wire N__22556;
    wire N__22555;
    wire N__22554;
    wire N__22553;
    wire N__22552;
    wire N__22551;
    wire N__22550;
    wire N__22549;
    wire N__22548;
    wire N__22543;
    wire N__22540;
    wire N__22539;
    wire N__22538;
    wire N__22535;
    wire N__22534;
    wire N__22533;
    wire N__22530;
    wire N__22529;
    wire N__22528;
    wire N__22525;
    wire N__22522;
    wire N__22519;
    wire N__22514;
    wire N__22509;
    wire N__22500;
    wire N__22487;
    wire N__22476;
    wire N__22473;
    wire N__22470;
    wire N__22467;
    wire N__22466;
    wire N__22463;
    wire N__22460;
    wire N__22455;
    wire N__22452;
    wire N__22451;
    wire N__22450;
    wire N__22447;
    wire N__22444;
    wire N__22441;
    wire N__22436;
    wire N__22433;
    wire N__22430;
    wire N__22427;
    wire N__22422;
    wire N__22419;
    wire N__22418;
    wire N__22415;
    wire N__22414;
    wire N__22411;
    wire N__22408;
    wire N__22405;
    wire N__22402;
    wire N__22395;
    wire N__22392;
    wire N__22389;
    wire N__22386;
    wire N__22385;
    wire N__22382;
    wire N__22379;
    wire N__22378;
    wire N__22375;
    wire N__22372;
    wire N__22369;
    wire N__22366;
    wire N__22359;
    wire N__22356;
    wire N__22353;
    wire N__22352;
    wire N__22351;
    wire N__22348;
    wire N__22345;
    wire N__22342;
    wire N__22339;
    wire N__22332;
    wire N__22331;
    wire N__22328;
    wire N__22325;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22315;
    wire N__22312;
    wire N__22309;
    wire N__22306;
    wire N__22303;
    wire N__22298;
    wire N__22293;
    wire N__22290;
    wire N__22289;
    wire N__22286;
    wire N__22283;
    wire N__22282;
    wire N__22279;
    wire N__22276;
    wire N__22273;
    wire N__22268;
    wire N__22263;
    wire N__22262;
    wire N__22259;
    wire N__22256;
    wire N__22253;
    wire N__22252;
    wire N__22249;
    wire N__22246;
    wire N__22243;
    wire N__22236;
    wire N__22233;
    wire N__22230;
    wire N__22227;
    wire N__22224;
    wire N__22221;
    wire N__22218;
    wire N__22215;
    wire N__22212;
    wire N__22209;
    wire N__22206;
    wire N__22203;
    wire N__22200;
    wire N__22197;
    wire N__22194;
    wire N__22193;
    wire N__22192;
    wire N__22191;
    wire N__22190;
    wire N__22189;
    wire N__22188;
    wire N__22187;
    wire N__22186;
    wire N__22185;
    wire N__22178;
    wire N__22175;
    wire N__22172;
    wire N__22171;
    wire N__22168;
    wire N__22165;
    wire N__22160;
    wire N__22159;
    wire N__22156;
    wire N__22151;
    wire N__22150;
    wire N__22147;
    wire N__22144;
    wire N__22143;
    wire N__22142;
    wire N__22141;
    wire N__22140;
    wire N__22139;
    wire N__22136;
    wire N__22131;
    wire N__22128;
    wire N__22123;
    wire N__22120;
    wire N__22117;
    wire N__22114;
    wire N__22111;
    wire N__22110;
    wire N__22109;
    wire N__22108;
    wire N__22107;
    wire N__22106;
    wire N__22105;
    wire N__22104;
    wire N__22103;
    wire N__22102;
    wire N__22101;
    wire N__22100;
    wire N__22099;
    wire N__22098;
    wire N__22089;
    wire N__22084;
    wire N__22077;
    wire N__22070;
    wire N__22059;
    wire N__22042;
    wire N__22029;
    wire N__22026;
    wire N__22023;
    wire N__22020;
    wire N__22019;
    wire N__22018;
    wire N__22017;
    wire N__22016;
    wire N__22015;
    wire N__22014;
    wire N__22013;
    wire N__22012;
    wire N__22009;
    wire N__22008;
    wire N__22005;
    wire N__22004;
    wire N__22003;
    wire N__22002;
    wire N__22001;
    wire N__22000;
    wire N__21997;
    wire N__21994;
    wire N__21991;
    wire N__21986;
    wire N__21985;
    wire N__21980;
    wire N__21977;
    wire N__21974;
    wire N__21971;
    wire N__21970;
    wire N__21969;
    wire N__21958;
    wire N__21949;
    wire N__21946;
    wire N__21941;
    wire N__21936;
    wire N__21935;
    wire N__21934;
    wire N__21933;
    wire N__21930;
    wire N__21929;
    wire N__21928;
    wire N__21927;
    wire N__21924;
    wire N__21923;
    wire N__21922;
    wire N__21921;
    wire N__21920;
    wire N__21919;
    wire N__21918;
    wire N__21917;
    wire N__21912;
    wire N__21905;
    wire N__21900;
    wire N__21897;
    wire N__21894;
    wire N__21881;
    wire N__21870;
    wire N__21855;
    wire N__21852;
    wire N__21849;
    wire N__21846;
    wire N__21845;
    wire N__21842;
    wire N__21839;
    wire N__21838;
    wire N__21835;
    wire N__21832;
    wire N__21829;
    wire N__21826;
    wire N__21823;
    wire N__21820;
    wire N__21813;
    wire N__21810;
    wire N__21807;
    wire N__21804;
    wire N__21803;
    wire N__21802;
    wire N__21801;
    wire N__21800;
    wire N__21799;
    wire N__21796;
    wire N__21795;
    wire N__21794;
    wire N__21793;
    wire N__21792;
    wire N__21791;
    wire N__21788;
    wire N__21787;
    wire N__21786;
    wire N__21783;
    wire N__21782;
    wire N__21781;
    wire N__21778;
    wire N__21777;
    wire N__21774;
    wire N__21771;
    wire N__21768;
    wire N__21765;
    wire N__21758;
    wire N__21755;
    wire N__21744;
    wire N__21733;
    wire N__21720;
    wire N__21719;
    wire N__21716;
    wire N__21713;
    wire N__21710;
    wire N__21707;
    wire N__21702;
    wire N__21699;
    wire N__21696;
    wire N__21693;
    wire N__21690;
    wire N__21687;
    wire N__21684;
    wire N__21681;
    wire N__21678;
    wire N__21675;
    wire N__21672;
    wire N__21669;
    wire N__21666;
    wire N__21663;
    wire N__21660;
    wire N__21657;
    wire N__21654;
    wire N__21651;
    wire N__21648;
    wire N__21645;
    wire N__21642;
    wire N__21639;
    wire N__21636;
    wire N__21633;
    wire N__21630;
    wire N__21627;
    wire N__21624;
    wire N__21621;
    wire N__21618;
    wire N__21615;
    wire N__21612;
    wire N__21609;
    wire N__21606;
    wire N__21603;
    wire N__21600;
    wire N__21597;
    wire N__21594;
    wire N__21591;
    wire N__21588;
    wire N__21585;
    wire N__21582;
    wire N__21579;
    wire N__21576;
    wire N__21573;
    wire N__21570;
    wire N__21567;
    wire N__21564;
    wire N__21561;
    wire N__21558;
    wire N__21555;
    wire N__21552;
    wire N__21549;
    wire N__21546;
    wire N__21543;
    wire N__21540;
    wire N__21537;
    wire N__21534;
    wire N__21531;
    wire N__21528;
    wire N__21525;
    wire N__21522;
    wire N__21519;
    wire N__21516;
    wire N__21513;
    wire N__21510;
    wire N__21507;
    wire N__21504;
    wire N__21501;
    wire N__21500;
    wire N__21497;
    wire N__21496;
    wire N__21493;
    wire N__21490;
    wire N__21487;
    wire N__21484;
    wire N__21477;
    wire N__21474;
    wire N__21471;
    wire N__21468;
    wire N__21465;
    wire N__21464;
    wire N__21461;
    wire N__21458;
    wire N__21455;
    wire N__21452;
    wire N__21451;
    wire N__21446;
    wire N__21443;
    wire N__21440;
    wire N__21435;
    wire N__21432;
    wire N__21429;
    wire N__21426;
    wire N__21423;
    wire N__21422;
    wire N__21421;
    wire N__21420;
    wire N__21417;
    wire N__21414;
    wire N__21413;
    wire N__21412;
    wire N__21407;
    wire N__21404;
    wire N__21401;
    wire N__21398;
    wire N__21395;
    wire N__21390;
    wire N__21381;
    wire N__21378;
    wire N__21375;
    wire N__21372;
    wire N__21369;
    wire N__21368;
    wire N__21365;
    wire N__21362;
    wire N__21357;
    wire N__21354;
    wire N__21351;
    wire N__21348;
    wire N__21345;
    wire N__21342;
    wire N__21339;
    wire N__21336;
    wire N__21333;
    wire N__21330;
    wire N__21327;
    wire N__21326;
    wire N__21323;
    wire N__21320;
    wire N__21317;
    wire N__21316;
    wire N__21313;
    wire N__21310;
    wire N__21307;
    wire N__21300;
    wire N__21297;
    wire N__21296;
    wire N__21295;
    wire N__21292;
    wire N__21289;
    wire N__21286;
    wire N__21283;
    wire N__21280;
    wire N__21277;
    wire N__21274;
    wire N__21271;
    wire N__21268;
    wire N__21261;
    wire N__21258;
    wire N__21255;
    wire N__21252;
    wire N__21249;
    wire N__21246;
    wire N__21245;
    wire N__21244;
    wire N__21241;
    wire N__21238;
    wire N__21235;
    wire N__21228;
    wire N__21227;
    wire N__21226;
    wire N__21223;
    wire N__21220;
    wire N__21217;
    wire N__21214;
    wire N__21207;
    wire N__21204;
    wire N__21201;
    wire N__21198;
    wire N__21195;
    wire N__21192;
    wire N__21189;
    wire N__21186;
    wire N__21183;
    wire N__21180;
    wire N__21177;
    wire N__21174;
    wire N__21171;
    wire N__21168;
    wire N__21165;
    wire N__21162;
    wire N__21159;
    wire N__21158;
    wire N__21155;
    wire N__21154;
    wire N__21151;
    wire N__21148;
    wire N__21145;
    wire N__21138;
    wire N__21135;
    wire N__21132;
    wire N__21129;
    wire N__21126;
    wire N__21123;
    wire N__21120;
    wire N__21117;
    wire N__21114;
    wire N__21111;
    wire N__21108;
    wire N__21105;
    wire N__21102;
    wire N__21099;
    wire N__21096;
    wire N__21093;
    wire N__21090;
    wire N__21089;
    wire N__21088;
    wire N__21085;
    wire N__21080;
    wire N__21075;
    wire N__21074;
    wire N__21073;
    wire N__21070;
    wire N__21067;
    wire N__21064;
    wire N__21061;
    wire N__21054;
    wire N__21051;
    wire N__21048;
    wire N__21045;
    wire N__21042;
    wire N__21041;
    wire N__21038;
    wire N__21037;
    wire N__21034;
    wire N__21029;
    wire N__21024;
    wire N__21023;
    wire N__21022;
    wire N__21019;
    wire N__21016;
    wire N__21013;
    wire N__21006;
    wire N__21003;
    wire N__21000;
    wire N__20997;
    wire N__20994;
    wire N__20991;
    wire N__20990;
    wire N__20989;
    wire N__20988;
    wire N__20983;
    wire N__20978;
    wire N__20973;
    wire N__20970;
    wire N__20969;
    wire N__20968;
    wire N__20967;
    wire N__20962;
    wire N__20957;
    wire N__20952;
    wire N__20951;
    wire N__20946;
    wire N__20943;
    wire N__20942;
    wire N__20941;
    wire N__20936;
    wire N__20933;
    wire N__20928;
    wire N__20925;
    wire N__20924;
    wire N__20923;
    wire N__20918;
    wire N__20915;
    wire N__20912;
    wire N__20907;
    wire N__20904;
    wire N__20901;
    wire N__20898;
    wire N__20895;
    wire N__20892;
    wire N__20889;
    wire N__20888;
    wire N__20885;
    wire N__20882;
    wire N__20877;
    wire N__20876;
    wire N__20875;
    wire N__20872;
    wire N__20869;
    wire N__20866;
    wire N__20863;
    wire N__20860;
    wire N__20857;
    wire N__20852;
    wire N__20849;
    wire N__20844;
    wire N__20841;
    wire N__20840;
    wire N__20837;
    wire N__20834;
    wire N__20831;
    wire N__20830;
    wire N__20825;
    wire N__20822;
    wire N__20817;
    wire N__20814;
    wire N__20811;
    wire N__20808;
    wire N__20805;
    wire N__20802;
    wire N__20799;
    wire N__20796;
    wire N__20793;
    wire N__20790;
    wire N__20787;
    wire N__20784;
    wire N__20781;
    wire N__20778;
    wire N__20775;
    wire N__20772;
    wire N__20769;
    wire N__20766;
    wire N__20763;
    wire N__20760;
    wire N__20757;
    wire N__20754;
    wire N__20751;
    wire N__20748;
    wire N__20745;
    wire N__20742;
    wire N__20739;
    wire N__20736;
    wire N__20733;
    wire N__20730;
    wire N__20727;
    wire N__20724;
    wire N__20721;
    wire N__20718;
    wire N__20715;
    wire N__20712;
    wire N__20709;
    wire N__20706;
    wire N__20703;
    wire N__20700;
    wire N__20697;
    wire N__20694;
    wire N__20691;
    wire N__20688;
    wire N__20685;
    wire N__20682;
    wire N__20679;
    wire N__20676;
    wire N__20673;
    wire N__20670;
    wire N__20667;
    wire N__20664;
    wire N__20661;
    wire N__20658;
    wire N__20655;
    wire N__20652;
    wire N__20649;
    wire N__20646;
    wire N__20643;
    wire N__20640;
    wire N__20637;
    wire N__20634;
    wire N__20631;
    wire N__20628;
    wire N__20625;
    wire N__20622;
    wire N__20619;
    wire N__20616;
    wire N__20613;
    wire N__20610;
    wire N__20607;
    wire N__20604;
    wire N__20601;
    wire N__20598;
    wire N__20595;
    wire N__20592;
    wire N__20589;
    wire N__20586;
    wire N__20583;
    wire N__20580;
    wire N__20577;
    wire N__20574;
    wire N__20571;
    wire N__20568;
    wire N__20565;
    wire N__20562;
    wire N__20559;
    wire N__20558;
    wire N__20555;
    wire N__20554;
    wire N__20551;
    wire N__20548;
    wire N__20545;
    wire N__20542;
    wire N__20539;
    wire N__20536;
    wire N__20533;
    wire N__20526;
    wire N__20523;
    wire N__20520;
    wire N__20517;
    wire N__20514;
    wire N__20511;
    wire N__20508;
    wire N__20505;
    wire N__20502;
    wire N__20499;
    wire N__20496;
    wire N__20493;
    wire N__20490;
    wire N__20487;
    wire N__20484;
    wire N__20481;
    wire N__20478;
    wire N__20475;
    wire N__20472;
    wire N__20469;
    wire N__20466;
    wire N__20463;
    wire N__20460;
    wire N__20457;
    wire N__20454;
    wire N__20451;
    wire N__20448;
    wire N__20445;
    wire N__20442;
    wire N__20439;
    wire N__20436;
    wire N__20433;
    wire N__20430;
    wire N__20427;
    wire N__20424;
    wire N__20421;
    wire N__20418;
    wire N__20415;
    wire N__20412;
    wire N__20409;
    wire N__20406;
    wire N__20403;
    wire N__20400;
    wire N__20397;
    wire N__20394;
    wire N__20391;
    wire N__20388;
    wire N__20385;
    wire N__20382;
    wire N__20379;
    wire N__20376;
    wire N__20373;
    wire N__20370;
    wire N__20367;
    wire N__20364;
    wire N__20361;
    wire N__20358;
    wire N__20355;
    wire N__20352;
    wire N__20351;
    wire N__20350;
    wire N__20347;
    wire N__20344;
    wire N__20341;
    wire N__20338;
    wire N__20331;
    wire N__20328;
    wire N__20327;
    wire N__20324;
    wire N__20323;
    wire N__20320;
    wire N__20317;
    wire N__20314;
    wire N__20307;
    wire N__20304;
    wire N__20301;
    wire N__20298;
    wire N__20295;
    wire N__20292;
    wire N__20289;
    wire N__20286;
    wire N__20283;
    wire N__20282;
    wire N__20279;
    wire N__20276;
    wire N__20273;
    wire N__20270;
    wire N__20267;
    wire N__20264;
    wire N__20263;
    wire N__20260;
    wire N__20257;
    wire N__20254;
    wire N__20247;
    wire N__20244;
    wire N__20241;
    wire N__20240;
    wire N__20235;
    wire N__20232;
    wire N__20231;
    wire N__20228;
    wire N__20225;
    wire N__20224;
    wire N__20217;
    wire N__20214;
    wire N__20211;
    wire N__20210;
    wire N__20209;
    wire N__20206;
    wire N__20203;
    wire N__20200;
    wire N__20197;
    wire N__20190;
    wire N__20187;
    wire N__20184;
    wire N__20181;
    wire N__20180;
    wire N__20179;
    wire N__20176;
    wire N__20173;
    wire N__20170;
    wire N__20167;
    wire N__20160;
    wire N__20157;
    wire N__20154;
    wire N__20151;
    wire N__20148;
    wire N__20145;
    wire N__20142;
    wire N__20139;
    wire N__20136;
    wire N__20133;
    wire N__20130;
    wire N__20127;
    wire N__20124;
    wire N__20121;
    wire N__20118;
    wire N__20115;
    wire N__20112;
    wire N__20109;
    wire N__20108;
    wire N__20105;
    wire N__20102;
    wire N__20101;
    wire N__20098;
    wire N__20095;
    wire N__20092;
    wire N__20087;
    wire N__20082;
    wire N__20079;
    wire N__20076;
    wire N__20073;
    wire N__20072;
    wire N__20069;
    wire N__20066;
    wire N__20065;
    wire N__20062;
    wire N__20059;
    wire N__20056;
    wire N__20049;
    wire N__20048;
    wire N__20047;
    wire N__20044;
    wire N__20041;
    wire N__20038;
    wire N__20035;
    wire N__20032;
    wire N__20029;
    wire N__20024;
    wire N__20019;
    wire N__20016;
    wire N__20013;
    wire N__20012;
    wire N__20009;
    wire N__20008;
    wire N__20005;
    wire N__20002;
    wire N__19999;
    wire N__19996;
    wire N__19993;
    wire N__19986;
    wire N__19983;
    wire N__19980;
    wire N__19977;
    wire N__19974;
    wire N__19973;
    wire N__19970;
    wire N__19967;
    wire N__19964;
    wire N__19961;
    wire N__19960;
    wire N__19957;
    wire N__19954;
    wire N__19951;
    wire N__19944;
    wire N__19941;
    wire N__19938;
    wire N__19935;
    wire N__19932;
    wire N__19929;
    wire N__19928;
    wire N__19925;
    wire N__19922;
    wire N__19921;
    wire N__19918;
    wire N__19915;
    wire N__19912;
    wire N__19905;
    wire N__19902;
    wire N__19899;
    wire N__19896;
    wire N__19893;
    wire N__19890;
    wire N__19887;
    wire N__19884;
    wire N__19881;
    wire N__19878;
    wire N__19875;
    wire N__19872;
    wire N__19869;
    wire N__19866;
    wire N__19863;
    wire N__19860;
    wire N__19857;
    wire N__19854;
    wire N__19851;
    wire N__19848;
    wire N__19845;
    wire N__19842;
    wire N__19839;
    wire N__19836;
    wire N__19833;
    wire N__19830;
    wire N__19827;
    wire N__19824;
    wire N__19821;
    wire N__19818;
    wire N__19815;
    wire N__19812;
    wire N__19809;
    wire N__19806;
    wire N__19803;
    wire N__19800;
    wire N__19797;
    wire N__19794;
    wire N__19791;
    wire N__19788;
    wire N__19785;
    wire N__19782;
    wire N__19779;
    wire N__19776;
    wire N__19773;
    wire N__19770;
    wire N__19767;
    wire N__19764;
    wire N__19761;
    wire N__19758;
    wire N__19755;
    wire N__19752;
    wire N__19749;
    wire N__19746;
    wire N__19743;
    wire N__19740;
    wire N__19737;
    wire N__19734;
    wire N__19731;
    wire N__19728;
    wire N__19725;
    wire N__19722;
    wire N__19719;
    wire N__19716;
    wire N__19713;
    wire N__19710;
    wire N__19707;
    wire N__19704;
    wire N__19701;
    wire N__19698;
    wire N__19695;
    wire N__19692;
    wire N__19689;
    wire N__19686;
    wire N__19683;
    wire N__19680;
    wire N__19677;
    wire N__19674;
    wire N__19671;
    wire N__19668;
    wire N__19665;
    wire N__19662;
    wire N__19659;
    wire N__19656;
    wire N__19653;
    wire N__19652;
    wire N__19651;
    wire N__19650;
    wire N__19649;
    wire N__19646;
    wire N__19643;
    wire N__19640;
    wire N__19639;
    wire N__19636;
    wire N__19635;
    wire N__19632;
    wire N__19627;
    wire N__19624;
    wire N__19621;
    wire N__19618;
    wire N__19615;
    wire N__19612;
    wire N__19609;
    wire N__19606;
    wire N__19603;
    wire N__19598;
    wire N__19597;
    wire N__19594;
    wire N__19587;
    wire N__19584;
    wire N__19581;
    wire N__19572;
    wire N__19571;
    wire N__19570;
    wire N__19569;
    wire N__19562;
    wire N__19559;
    wire N__19554;
    wire N__19553;
    wire N__19552;
    wire N__19551;
    wire N__19542;
    wire N__19539;
    wire N__19538;
    wire N__19535;
    wire N__19532;
    wire N__19529;
    wire N__19524;
    wire N__19523;
    wire N__19520;
    wire N__19519;
    wire N__19516;
    wire N__19513;
    wire N__19510;
    wire N__19503;
    wire N__19502;
    wire N__19501;
    wire N__19498;
    wire N__19495;
    wire N__19492;
    wire N__19489;
    wire N__19482;
    wire N__19479;
    wire N__19476;
    wire N__19473;
    wire N__19470;
    wire N__19467;
    wire N__19464;
    wire N__19461;
    wire N__19458;
    wire N__19455;
    wire N__19454;
    wire N__19453;
    wire N__19452;
    wire N__19451;
    wire N__19450;
    wire N__19447;
    wire N__19442;
    wire N__19439;
    wire N__19436;
    wire N__19433;
    wire N__19430;
    wire N__19419;
    wire N__19416;
    wire N__19415;
    wire N__19414;
    wire N__19411;
    wire N__19408;
    wire N__19405;
    wire N__19402;
    wire N__19395;
    wire N__19394;
    wire N__19393;
    wire N__19390;
    wire N__19387;
    wire N__19384;
    wire N__19381;
    wire N__19378;
    wire N__19371;
    wire N__19370;
    wire N__19369;
    wire N__19366;
    wire N__19363;
    wire N__19360;
    wire N__19357;
    wire N__19354;
    wire N__19347;
    wire N__19346;
    wire N__19345;
    wire N__19342;
    wire N__19339;
    wire N__19336;
    wire N__19333;
    wire N__19330;
    wire N__19323;
    wire N__19320;
    wire N__19317;
    wire N__19316;
    wire N__19315;
    wire N__19312;
    wire N__19309;
    wire N__19306;
    wire N__19299;
    wire N__19298;
    wire N__19297;
    wire N__19294;
    wire N__19291;
    wire N__19288;
    wire N__19285;
    wire N__19278;
    wire N__19275;
    wire N__19272;
    wire N__19269;
    wire N__19266;
    wire N__19263;
    wire N__19260;
    wire N__19257;
    wire N__19256;
    wire N__19255;
    wire N__19252;
    wire N__19249;
    wire N__19246;
    wire N__19239;
    wire N__19238;
    wire N__19237;
    wire N__19234;
    wire N__19231;
    wire N__19228;
    wire N__19221;
    wire N__19220;
    wire N__19219;
    wire N__19216;
    wire N__19213;
    wire N__19210;
    wire N__19203;
    wire N__19200;
    wire N__19199;
    wire N__19198;
    wire N__19195;
    wire N__19190;
    wire N__19185;
    wire N__19182;
    wire N__19179;
    wire N__19176;
    wire N__19173;
    wire N__19172;
    wire N__19171;
    wire N__19168;
    wire N__19163;
    wire N__19158;
    wire N__19155;
    wire N__19152;
    wire N__19149;
    wire N__19146;
    wire N__19143;
    wire N__19140;
    wire N__19137;
    wire N__19134;
    wire N__19131;
    wire N__19128;
    wire N__19125;
    wire N__19122;
    wire N__19119;
    wire N__19116;
    wire N__19113;
    wire N__19110;
    wire N__19107;
    wire N__19104;
    wire N__19101;
    wire N__19098;
    wire N__19095;
    wire N__19092;
    wire N__19089;
    wire N__19088;
    wire N__19085;
    wire N__19082;
    wire N__19077;
    wire N__19074;
    wire N__19071;
    wire N__19068;
    wire N__19067;
    wire N__19066;
    wire N__19063;
    wire N__19058;
    wire N__19053;
    wire N__19050;
    wire N__19047;
    wire N__19044;
    wire N__19041;
    wire N__19040;
    wire N__19039;
    wire N__19036;
    wire N__19035;
    wire N__19034;
    wire N__19031;
    wire N__19030;
    wire N__19029;
    wire N__19028;
    wire N__19027;
    wire N__19026;
    wire N__19025;
    wire N__19024;
    wire N__19023;
    wire N__19022;
    wire N__19015;
    wire N__19008;
    wire N__19001;
    wire N__18994;
    wire N__18989;
    wire N__18978;
    wire N__18977;
    wire N__18976;
    wire N__18975;
    wire N__18974;
    wire N__18973;
    wire N__18972;
    wire N__18971;
    wire N__18968;
    wire N__18965;
    wire N__18964;
    wire N__18961;
    wire N__18958;
    wire N__18955;
    wire N__18954;
    wire N__18951;
    wire N__18950;
    wire N__18949;
    wire N__18948;
    wire N__18947;
    wire N__18946;
    wire N__18945;
    wire N__18942;
    wire N__18939;
    wire N__18936;
    wire N__18931;
    wire N__18928;
    wire N__18925;
    wire N__18914;
    wire N__18901;
    wire N__18888;
    wire N__18885;
    wire N__18882;
    wire N__18879;
    wire N__18876;
    wire N__18873;
    wire N__18870;
    wire N__18867;
    wire N__18864;
    wire N__18863;
    wire N__18860;
    wire N__18857;
    wire N__18852;
    wire N__18849;
    wire N__18846;
    wire N__18843;
    wire N__18840;
    wire N__18837;
    wire N__18834;
    wire N__18831;
    wire N__18828;
    wire N__18825;
    wire N__18822;
    wire N__18819;
    wire N__18816;
    wire N__18813;
    wire N__18810;
    wire N__18807;
    wire N__18804;
    wire N__18801;
    wire N__18798;
    wire N__18795;
    wire N__18792;
    wire N__18789;
    wire N__18786;
    wire N__18783;
    wire N__18780;
    wire N__18777;
    wire N__18774;
    wire N__18771;
    wire N__18768;
    wire N__18765;
    wire N__18762;
    wire N__18759;
    wire N__18756;
    wire N__18753;
    wire N__18750;
    wire N__18747;
    wire N__18744;
    wire N__18741;
    wire N__18738;
    wire N__18735;
    wire N__18732;
    wire N__18729;
    wire N__18726;
    wire N__18723;
    wire N__18720;
    wire N__18717;
    wire N__18714;
    wire N__18711;
    wire N__18708;
    wire N__18705;
    wire N__18702;
    wire N__18699;
    wire N__18696;
    wire N__18693;
    wire N__18690;
    wire N__18687;
    wire N__18684;
    wire N__18681;
    wire N__18678;
    wire N__18675;
    wire N__18672;
    wire N__18669;
    wire N__18666;
    wire N__18663;
    wire N__18660;
    wire N__18657;
    wire N__18654;
    wire N__18651;
    wire N__18648;
    wire N__18645;
    wire N__18642;
    wire N__18639;
    wire N__18636;
    wire N__18633;
    wire N__18630;
    wire N__18627;
    wire N__18624;
    wire N__18621;
    wire N__18618;
    wire N__18615;
    wire N__18612;
    wire N__18609;
    wire N__18606;
    wire N__18603;
    wire N__18600;
    wire N__18597;
    wire N__18594;
    wire N__18591;
    wire N__18588;
    wire N__18585;
    wire N__18582;
    wire N__18579;
    wire N__18576;
    wire N__18573;
    wire N__18570;
    wire N__18567;
    wire N__18564;
    wire N__18561;
    wire N__18558;
    wire N__18555;
    wire N__18552;
    wire N__18549;
    wire N__18546;
    wire N__18543;
    wire N__18540;
    wire N__18537;
    wire N__18534;
    wire N__18531;
    wire N__18530;
    wire N__18529;
    wire N__18526;
    wire N__18523;
    wire N__18520;
    wire N__18519;
    wire N__18518;
    wire N__18517;
    wire N__18516;
    wire N__18515;
    wire N__18508;
    wire N__18507;
    wire N__18506;
    wire N__18505;
    wire N__18504;
    wire N__18503;
    wire N__18500;
    wire N__18499;
    wire N__18496;
    wire N__18493;
    wire N__18492;
    wire N__18491;
    wire N__18488;
    wire N__18485;
    wire N__18482;
    wire N__18473;
    wire N__18456;
    wire N__18447;
    wire N__18446;
    wire N__18443;
    wire N__18440;
    wire N__18435;
    wire N__18434;
    wire N__18433;
    wire N__18430;
    wire N__18427;
    wire N__18424;
    wire N__18417;
    wire N__18414;
    wire N__18411;
    wire N__18408;
    wire N__18407;
    wire N__18404;
    wire N__18401;
    wire N__18396;
    wire N__18393;
    wire N__18392;
    wire N__18389;
    wire N__18388;
    wire N__18387;
    wire N__18384;
    wire N__18383;
    wire N__18382;
    wire N__18381;
    wire N__18380;
    wire N__18379;
    wire N__18370;
    wire N__18369;
    wire N__18368;
    wire N__18365;
    wire N__18364;
    wire N__18361;
    wire N__18360;
    wire N__18359;
    wire N__18358;
    wire N__18355;
    wire N__18352;
    wire N__18351;
    wire N__18348;
    wire N__18345;
    wire N__18342;
    wire N__18331;
    wire N__18318;
    wire N__18309;
    wire N__18306;
    wire N__18303;
    wire N__18300;
    wire N__18297;
    wire N__18294;
    wire N__18291;
    wire N__18288;
    wire N__18285;
    wire N__18282;
    wire N__18279;
    wire N__18276;
    wire N__18273;
    wire N__18270;
    wire N__18267;
    wire N__18264;
    wire N__18261;
    wire N__18258;
    wire N__18255;
    wire N__18252;
    wire N__18249;
    wire N__18248;
    wire N__18245;
    wire N__18242;
    wire N__18239;
    wire N__18236;
    wire N__18235;
    wire N__18234;
    wire N__18233;
    wire N__18228;
    wire N__18225;
    wire N__18222;
    wire N__18219;
    wire N__18210;
    wire N__18207;
    wire N__18204;
    wire N__18201;
    wire N__18198;
    wire N__18195;
    wire N__18192;
    wire N__18189;
    wire N__18186;
    wire N__18183;
    wire N__18180;
    wire N__18177;
    wire N__18174;
    wire N__18173;
    wire N__18172;
    wire N__18169;
    wire N__18166;
    wire N__18163;
    wire N__18158;
    wire N__18153;
    wire N__18150;
    wire N__18147;
    wire N__18144;
    wire N__18141;
    wire N__18140;
    wire N__18137;
    wire N__18134;
    wire N__18133;
    wire N__18130;
    wire N__18127;
    wire N__18124;
    wire N__18121;
    wire N__18118;
    wire N__18111;
    wire N__18110;
    wire N__18107;
    wire N__18104;
    wire N__18101;
    wire N__18100;
    wire N__18097;
    wire N__18094;
    wire N__18091;
    wire N__18088;
    wire N__18085;
    wire N__18078;
    wire N__18077;
    wire N__18074;
    wire N__18071;
    wire N__18068;
    wire N__18067;
    wire N__18064;
    wire N__18061;
    wire N__18058;
    wire N__18055;
    wire N__18052;
    wire N__18045;
    wire N__18042;
    wire N__18039;
    wire N__18036;
    wire N__18035;
    wire N__18034;
    wire N__18029;
    wire N__18026;
    wire N__18023;
    wire N__18018;
    wire N__18015;
    wire N__18012;
    wire N__18011;
    wire N__18008;
    wire N__18007;
    wire N__18004;
    wire N__18001;
    wire N__17998;
    wire N__17993;
    wire N__17988;
    wire N__17985;
    wire N__17982;
    wire N__17979;
    wire N__17976;
    wire N__17973;
    wire N__17970;
    wire N__17967;
    wire N__17966;
    wire N__17963;
    wire N__17962;
    wire N__17959;
    wire N__17954;
    wire N__17949;
    wire N__17946;
    wire N__17943;
    wire N__17942;
    wire N__17941;
    wire N__17938;
    wire N__17935;
    wire N__17932;
    wire N__17929;
    wire N__17926;
    wire N__17919;
    wire N__17916;
    wire N__17913;
    wire N__17910;
    wire N__17907;
    wire N__17904;
    wire N__17901;
    wire N__17898;
    wire N__17895;
    wire N__17892;
    wire N__17889;
    wire N__17886;
    wire N__17883;
    wire N__17880;
    wire N__17877;
    wire N__17874;
    wire N__17871;
    wire N__17868;
    wire N__17865;
    wire N__17862;
    wire N__17859;
    wire N__17856;
    wire N__17855;
    wire N__17854;
    wire N__17851;
    wire N__17846;
    wire N__17841;
    wire N__17838;
    wire N__17835;
    wire N__17832;
    wire N__17829;
    wire N__17826;
    wire N__17823;
    wire N__17822;
    wire N__17817;
    wire N__17814;
    wire N__17813;
    wire N__17808;
    wire N__17807;
    wire N__17804;
    wire N__17801;
    wire N__17798;
    wire N__17795;
    wire N__17792;
    wire N__17789;
    wire N__17784;
    wire N__17781;
    wire N__17778;
    wire N__17775;
    wire N__17772;
    wire N__17769;
    wire N__17766;
    wire N__17763;
    wire N__17760;
    wire N__17757;
    wire N__17754;
    wire N__17751;
    wire N__17748;
    wire N__17745;
    wire N__17742;
    wire N__17739;
    wire N__17736;
    wire N__17733;
    wire N__17730;
    wire N__17727;
    wire N__17724;
    wire N__17721;
    wire N__17718;
    wire N__17715;
    wire N__17712;
    wire N__17709;
    wire N__17706;
    wire N__17703;
    wire N__17700;
    wire N__17697;
    wire N__17694;
    wire N__17691;
    wire N__17688;
    wire N__17685;
    wire N__17682;
    wire N__17679;
    wire N__17676;
    wire N__17673;
    wire N__17670;
    wire N__17667;
    wire N__17664;
    wire N__17661;
    wire N__17658;
    wire N__17655;
    wire N__17652;
    wire N__17649;
    wire N__17646;
    wire N__17643;
    wire N__17640;
    wire N__17637;
    wire N__17634;
    wire N__17631;
    wire N__17628;
    wire N__17625;
    wire N__17622;
    wire N__17619;
    wire N__17616;
    wire N__17613;
    wire N__17610;
    wire N__17607;
    wire N__17604;
    wire N__17601;
    wire N__17598;
    wire N__17595;
    wire N__17594;
    wire N__17593;
    wire N__17592;
    wire N__17591;
    wire N__17590;
    wire N__17589;
    wire N__17588;
    wire N__17585;
    wire N__17584;
    wire N__17581;
    wire N__17578;
    wire N__17577;
    wire N__17576;
    wire N__17573;
    wire N__17572;
    wire N__17569;
    wire N__17568;
    wire N__17565;
    wire N__17562;
    wire N__17561;
    wire N__17558;
    wire N__17555;
    wire N__17546;
    wire N__17529;
    wire N__17520;
    wire N__17517;
    wire N__17514;
    wire N__17511;
    wire N__17508;
    wire N__17505;
    wire N__17504;
    wire N__17503;
    wire N__17502;
    wire N__17501;
    wire N__17500;
    wire N__17499;
    wire N__17490;
    wire N__17487;
    wire N__17486;
    wire N__17483;
    wire N__17482;
    wire N__17479;
    wire N__17478;
    wire N__17477;
    wire N__17476;
    wire N__17475;
    wire N__17474;
    wire N__17471;
    wire N__17466;
    wire N__17457;
    wire N__17448;
    wire N__17439;
    wire N__17436;
    wire N__17433;
    wire N__17430;
    wire N__17427;
    wire N__17424;
    wire N__17421;
    wire N__17418;
    wire N__17415;
    wire N__17412;
    wire N__17409;
    wire N__17406;
    wire N__17403;
    wire N__17400;
    wire N__17397;
    wire N__17394;
    wire N__17391;
    wire N__17388;
    wire N__17385;
    wire N__17382;
    wire N__17379;
    wire N__17376;
    wire N__17373;
    wire N__17370;
    wire N__17367;
    wire N__17364;
    wire N__17361;
    wire N__17358;
    wire N__17355;
    wire N__17352;
    wire N__17349;
    wire N__17346;
    wire N__17343;
    wire N__17340;
    wire N__17337;
    wire N__17334;
    wire N__17331;
    wire N__17328;
    wire N__17325;
    wire N__17322;
    wire N__17319;
    wire N__17316;
    wire N__17313;
    wire N__17310;
    wire N__17307;
    wire N__17304;
    wire N__17301;
    wire N__17298;
    wire N__17295;
    wire N__17292;
    wire N__17291;
    wire N__17290;
    wire N__17289;
    wire N__17288;
    wire N__17285;
    wire N__17284;
    wire N__17281;
    wire N__17278;
    wire N__17273;
    wire N__17270;
    wire N__17267;
    wire N__17260;
    wire N__17253;
    wire N__17250;
    wire N__17247;
    wire N__17244;
    wire N__17243;
    wire N__17240;
    wire N__17237;
    wire N__17232;
    wire N__17229;
    wire N__17226;
    wire N__17223;
    wire N__17220;
    wire N__17217;
    wire N__17214;
    wire N__17211;
    wire N__17208;
    wire N__17205;
    wire N__17202;
    wire N__17199;
    wire N__17198;
    wire N__17195;
    wire N__17194;
    wire N__17191;
    wire N__17188;
    wire N__17185;
    wire N__17178;
    wire N__17175;
    wire N__17172;
    wire N__17171;
    wire N__17170;
    wire N__17167;
    wire N__17164;
    wire N__17161;
    wire N__17156;
    wire N__17151;
    wire N__17148;
    wire N__17147;
    wire N__17146;
    wire N__17143;
    wire N__17140;
    wire N__17137;
    wire N__17134;
    wire N__17131;
    wire N__17124;
    wire N__17121;
    wire N__17118;
    wire N__17115;
    wire N__17112;
    wire N__17111;
    wire N__17110;
    wire N__17107;
    wire N__17104;
    wire N__17101;
    wire N__17098;
    wire N__17095;
    wire N__17088;
    wire N__17087;
    wire N__17084;
    wire N__17081;
    wire N__17080;
    wire N__17077;
    wire N__17074;
    wire N__17071;
    wire N__17068;
    wire N__17065;
    wire N__17058;
    wire N__17055;
    wire N__17052;
    wire N__17049;
    wire N__17046;
    wire N__17043;
    wire N__17040;
    wire N__17037;
    wire N__17034;
    wire N__17031;
    wire N__17028;
    wire N__17027;
    wire N__17026;
    wire N__17023;
    wire N__17020;
    wire N__17017;
    wire N__17014;
    wire N__17011;
    wire N__17004;
    wire N__17003;
    wire N__17002;
    wire N__17001;
    wire N__17000;
    wire N__16999;
    wire N__16996;
    wire N__16991;
    wire N__16988;
    wire N__16985;
    wire N__16982;
    wire N__16973;
    wire N__16970;
    wire N__16967;
    wire N__16962;
    wire N__16959;
    wire N__16956;
    wire N__16953;
    wire N__16950;
    wire N__16947;
    wire N__16944;
    wire N__16941;
    wire N__16938;
    wire N__16935;
    wire N__16932;
    wire N__16929;
    wire N__16926;
    wire N__16923;
    wire N__16920;
    wire N__16917;
    wire N__16914;
    wire N__16911;
    wire N__16908;
    wire N__16905;
    wire N__16904;
    wire N__16901;
    wire N__16900;
    wire N__16897;
    wire N__16894;
    wire N__16891;
    wire N__16886;
    wire N__16881;
    wire N__16878;
    wire N__16875;
    wire N__16874;
    wire N__16869;
    wire N__16866;
    wire N__16865;
    wire N__16862;
    wire N__16859;
    wire N__16854;
    wire N__16853;
    wire N__16850;
    wire N__16847;
    wire N__16842;
    wire N__16841;
    wire N__16836;
    wire N__16833;
    wire N__16830;
    wire N__16827;
    wire N__16826;
    wire N__16825;
    wire N__16824;
    wire N__16823;
    wire N__16822;
    wire N__16819;
    wire N__16816;
    wire N__16813;
    wire N__16810;
    wire N__16807;
    wire N__16804;
    wire N__16803;
    wire N__16800;
    wire N__16795;
    wire N__16792;
    wire N__16789;
    wire N__16786;
    wire N__16783;
    wire N__16778;
    wire N__16775;
    wire N__16768;
    wire N__16765;
    wire N__16760;
    wire N__16755;
    wire N__16754;
    wire N__16753;
    wire N__16746;
    wire N__16743;
    wire N__16742;
    wire N__16739;
    wire N__16736;
    wire N__16735;
    wire N__16734;
    wire N__16725;
    wire N__16722;
    wire N__16721;
    wire N__16720;
    wire N__16719;
    wire N__16710;
    wire N__16707;
    wire N__16704;
    wire N__16703;
    wire N__16702;
    wire N__16697;
    wire N__16694;
    wire N__16691;
    wire N__16686;
    wire N__16683;
    wire N__16682;
    wire N__16679;
    wire N__16678;
    wire N__16675;
    wire N__16672;
    wire N__16669;
    wire N__16664;
    wire N__16659;
    wire N__16656;
    wire N__16655;
    wire N__16652;
    wire N__16649;
    wire N__16648;
    wire N__16645;
    wire N__16642;
    wire N__16639;
    wire N__16636;
    wire N__16633;
    wire N__16626;
    wire N__16623;
    wire N__16620;
    wire N__16619;
    wire N__16618;
    wire N__16615;
    wire N__16612;
    wire N__16609;
    wire N__16604;
    wire N__16599;
    wire N__16596;
    wire N__16595;
    wire N__16592;
    wire N__16589;
    wire N__16586;
    wire N__16581;
    wire N__16580;
    wire N__16577;
    wire N__16574;
    wire N__16569;
    wire N__16566;
    wire N__16563;
    wire N__16560;
    wire N__16557;
    wire N__16554;
    wire N__16551;
    wire N__16548;
    wire N__16545;
    wire N__16542;
    wire N__16539;
    wire N__16536;
    wire N__16533;
    wire N__16530;
    wire N__16527;
    wire N__16524;
    wire N__16523;
    wire N__16522;
    wire N__16521;
    wire N__16518;
    wire N__16515;
    wire N__16514;
    wire N__16513;
    wire N__16512;
    wire N__16511;
    wire N__16510;
    wire N__16509;
    wire N__16508;
    wire N__16507;
    wire N__16506;
    wire N__16505;
    wire N__16502;
    wire N__16495;
    wire N__16484;
    wire N__16473;
    wire N__16464;
    wire N__16463;
    wire N__16462;
    wire N__16459;
    wire N__16454;
    wire N__16449;
    wire N__16446;
    wire N__16443;
    wire N__16440;
    wire N__16437;
    wire N__16434;
    wire N__16431;
    wire N__16428;
    wire N__16425;
    wire N__16422;
    wire N__16419;
    wire N__16416;
    wire N__16413;
    wire N__16410;
    wire N__16407;
    wire N__16404;
    wire N__16401;
    wire N__16398;
    wire N__16395;
    wire N__16392;
    wire N__16389;
    wire N__16386;
    wire N__16385;
    wire N__16382;
    wire N__16379;
    wire N__16374;
    wire N__16371;
    wire N__16368;
    wire N__16365;
    wire N__16362;
    wire N__16359;
    wire N__16356;
    wire N__16353;
    wire N__16350;
    wire N__16349;
    wire N__16348;
    wire N__16345;
    wire N__16342;
    wire N__16339;
    wire N__16336;
    wire N__16333;
    wire N__16326;
    wire N__16323;
    wire N__16322;
    wire N__16319;
    wire N__16318;
    wire N__16315;
    wire N__16312;
    wire N__16309;
    wire N__16302;
    wire N__16299;
    wire N__16296;
    wire N__16295;
    wire N__16294;
    wire N__16291;
    wire N__16288;
    wire N__16285;
    wire N__16280;
    wire N__16275;
    wire N__16272;
    wire N__16271;
    wire N__16268;
    wire N__16267;
    wire N__16264;
    wire N__16261;
    wire N__16258;
    wire N__16251;
    wire N__16248;
    wire N__16245;
    wire N__16242;
    wire N__16241;
    wire N__16240;
    wire N__16237;
    wire N__16234;
    wire N__16229;
    wire N__16224;
    wire N__16221;
    wire N__16220;
    wire N__16219;
    wire N__16216;
    wire N__16211;
    wire N__16206;
    wire N__16203;
    wire N__16202;
    wire N__16201;
    wire N__16198;
    wire N__16195;
    wire N__16190;
    wire N__16185;
    wire N__16182;
    wire N__16179;
    wire N__16178;
    wire N__16173;
    wire N__16172;
    wire N__16169;
    wire N__16166;
    wire N__16163;
    wire N__16158;
    wire N__16155;
    wire N__16152;
    wire N__16151;
    wire N__16150;
    wire N__16147;
    wire N__16144;
    wire N__16141;
    wire N__16134;
    wire N__16131;
    wire N__16130;
    wire N__16129;
    wire N__16126;
    wire N__16123;
    wire N__16120;
    wire N__16117;
    wire N__16110;
    wire N__16107;
    wire N__16104;
    wire N__16103;
    wire N__16102;
    wire N__16099;
    wire N__16096;
    wire N__16093;
    wire N__16090;
    wire N__16083;
    wire N__16080;
    wire N__16077;
    wire N__16074;
    wire N__16071;
    wire N__16068;
    wire N__16065;
    wire N__16062;
    wire N__16061;
    wire N__16060;
    wire N__16055;
    wire N__16052;
    wire N__16049;
    wire N__16044;
    wire N__16043;
    wire N__16042;
    wire N__16037;
    wire N__16034;
    wire N__16031;
    wire N__16026;
    wire N__16023;
    wire N__16022;
    wire N__16021;
    wire N__16018;
    wire N__16013;
    wire N__16008;
    wire N__16005;
    wire N__16004;
    wire N__16003;
    wire N__15998;
    wire N__15995;
    wire N__15992;
    wire N__15987;
    wire N__15984;
    wire N__15983;
    wire N__15980;
    wire N__15979;
    wire N__15974;
    wire N__15971;
    wire N__15968;
    wire N__15963;
    wire N__15960;
    wire N__15959;
    wire N__15958;
    wire N__15953;
    wire N__15950;
    wire N__15947;
    wire N__15942;
    wire N__15939;
    wire N__15938;
    wire N__15935;
    wire N__15934;
    wire N__15929;
    wire N__15926;
    wire N__15923;
    wire N__15918;
    wire N__15915;
    wire N__15912;
    wire N__15909;
    wire N__15906;
    wire N__15903;
    wire N__15900;
    wire N__15899;
    wire N__15894;
    wire N__15891;
    wire N__15888;
    wire N__15887;
    wire N__15886;
    wire N__15883;
    wire N__15882;
    wire N__15873;
    wire N__15870;
    wire N__15869;
    wire N__15868;
    wire N__15867;
    wire N__15858;
    wire N__15855;
    wire N__15852;
    wire N__15849;
    wire N__15846;
    wire N__15843;
    wire N__15840;
    wire N__15837;
    wire N__15834;
    wire N__15831;
    wire N__15830;
    wire N__15827;
    wire N__15824;
    wire N__15821;
    wire N__15816;
    wire N__15813;
    wire N__15810;
    wire N__15807;
    wire N__15804;
    wire N__15801;
    wire N__15798;
    wire N__15795;
    wire N__15792;
    wire N__15789;
    wire N__15786;
    wire N__15783;
    wire N__15780;
    wire N__15777;
    wire N__15774;
    wire N__15771;
    wire N__15768;
    wire N__15765;
    wire N__15762;
    wire N__15759;
    wire N__15756;
    wire N__15753;
    wire N__15750;
    wire N__15747;
    wire N__15744;
    wire N__15741;
    wire N__15738;
    wire N__15735;
    wire N__15732;
    wire N__15729;
    wire N__15726;
    wire N__15725;
    wire N__15722;
    wire N__15719;
    wire N__15714;
    wire N__15711;
    wire N__15708;
    wire N__15705;
    wire N__15704;
    wire N__15701;
    wire N__15698;
    wire N__15693;
    wire N__15692;
    wire N__15687;
    wire N__15684;
    wire N__15681;
    wire N__15678;
    wire N__15675;
    wire N__15672;
    wire N__15669;
    wire N__15666;
    wire N__15663;
    wire N__15660;
    wire N__15657;
    wire N__15654;
    wire N__15651;
    wire N__15648;
    wire N__15645;
    wire N__15642;
    wire N__15639;
    wire N__15636;
    wire N__15633;
    wire N__15630;
    wire N__15627;
    wire N__15624;
    wire N__15621;
    wire N__15618;
    wire N__15615;
    wire N__15612;
    wire N__15609;
    wire N__15606;
    wire N__15603;
    wire N__15600;
    wire N__15597;
    wire N__15594;
    wire N__15591;
    wire N__15588;
    wire N__15585;
    wire N__15582;
    wire N__15579;
    wire N__15576;
    wire N__15575;
    wire N__15574;
    wire N__15571;
    wire N__15568;
    wire N__15565;
    wire N__15560;
    wire N__15555;
    wire N__15552;
    wire N__15549;
    wire N__15546;
    wire N__15543;
    wire N__15540;
    wire N__15537;
    wire N__15534;
    wire N__15531;
    wire N__15528;
    wire N__15525;
    wire N__15522;
    wire N__15519;
    wire N__15516;
    wire N__15513;
    wire N__15510;
    wire N__15507;
    wire N__15504;
    wire N__15501;
    wire N__15498;
    wire N__15495;
    wire N__15492;
    wire N__15489;
    wire N__15486;
    wire N__15483;
    wire N__15480;
    wire N__15477;
    wire N__15474;
    wire N__15471;
    wire N__15468;
    wire N__15465;
    wire N__15462;
    wire N__15459;
    wire N__15456;
    wire N__15453;
    wire N__15450;
    wire N__15447;
    wire N__15444;
    wire N__15441;
    wire N__15438;
    wire N__15435;
    wire N__15432;
    wire N__15429;
    wire N__15426;
    wire N__15423;
    wire N__15420;
    wire N__15417;
    wire N__15414;
    wire N__15411;
    wire N__15408;
    wire N__15405;
    wire N__15402;
    wire N__15399;
    wire N__15396;
    wire N__15393;
    wire N__15390;
    wire N__15387;
    wire N__15384;
    wire N__15381;
    wire N__15378;
    wire N__15375;
    wire N__15372;
    wire N__15369;
    wire N__15366;
    wire N__15363;
    wire N__15360;
    wire N__15357;
    wire N__15354;
    wire N__15351;
    wire N__15348;
    wire N__15345;
    wire N__15342;
    wire N__15339;
    wire N__15336;
    wire N__15333;
    wire N__15330;
    wire N__15327;
    wire N__15324;
    wire N__15321;
    wire N__15318;
    wire N__15315;
    wire N__15312;
    wire N__15309;
    wire N__15306;
    wire N__15303;
    wire N__15300;
    wire N__15297;
    wire N__15294;
    wire N__15291;
    wire N__15288;
    wire N__15285;
    wire N__15282;
    wire N__15279;
    wire N__15276;
    wire N__15275;
    wire N__15272;
    wire N__15271;
    wire N__15270;
    wire N__15267;
    wire N__15266;
    wire N__15263;
    wire N__15260;
    wire N__15257;
    wire N__15254;
    wire N__15251;
    wire N__15246;
    wire N__15243;
    wire N__15240;
    wire N__15237;
    wire N__15232;
    wire N__15229;
    wire N__15226;
    wire N__15219;
    wire N__15216;
    wire N__15213;
    wire N__15210;
    wire N__15207;
    wire N__15204;
    wire N__15201;
    wire N__15198;
    wire N__15195;
    wire N__15192;
    wire N__15189;
    wire N__15186;
    wire N__15183;
    wire N__15180;
    wire N__15177;
    wire N__15174;
    wire N__15171;
    wire N__15168;
    wire N__15165;
    wire N__15162;
    wire N__15159;
    wire N__15156;
    wire N__15153;
    wire N__15150;
    wire N__15147;
    wire N__15144;
    wire N__15141;
    wire N__15138;
    wire N__15135;
    wire N__15132;
    wire N__15129;
    wire N__15126;
    wire N__15123;
    wire N__15120;
    wire N__15119;
    wire N__15118;
    wire N__15115;
    wire N__15112;
    wire N__15109;
    wire N__15106;
    wire N__15103;
    wire N__15096;
    wire N__15095;
    wire N__15092;
    wire N__15089;
    wire N__15088;
    wire N__15085;
    wire N__15082;
    wire N__15079;
    wire N__15074;
    wire N__15069;
    wire N__15066;
    wire N__15063;
    wire N__15060;
    wire N__15057;
    wire N__15056;
    wire N__15055;
    wire N__15052;
    wire N__15049;
    wire N__15046;
    wire N__15043;
    wire N__15036;
    wire N__15033;
    wire N__15030;
    wire N__15029;
    wire N__15028;
    wire N__15025;
    wire N__15022;
    wire N__15019;
    wire N__15016;
    wire N__15009;
    wire N__15006;
    wire N__15003;
    wire N__15000;
    wire N__14999;
    wire N__14998;
    wire N__14995;
    wire N__14992;
    wire N__14989;
    wire N__14986;
    wire N__14979;
    wire N__14976;
    wire N__14975;
    wire N__14972;
    wire N__14971;
    wire N__14968;
    wire N__14965;
    wire N__14962;
    wire N__14955;
    wire N__14952;
    wire N__14949;
    wire N__14946;
    wire N__14943;
    wire N__14940;
    wire N__14939;
    wire N__14938;
    wire N__14935;
    wire N__14930;
    wire N__14929;
    wire N__14928;
    wire N__14927;
    wire N__14924;
    wire N__14921;
    wire N__14918;
    wire N__14915;
    wire N__14912;
    wire N__14909;
    wire N__14898;
    wire N__14895;
    wire N__14892;
    wire N__14889;
    wire N__14886;
    wire N__14883;
    wire N__14882;
    wire N__14879;
    wire N__14876;
    wire N__14871;
    wire N__14870;
    wire N__14865;
    wire N__14862;
    wire N__14859;
    wire N__14856;
    wire N__14853;
    wire N__14850;
    wire N__14847;
    wire N__14844;
    wire N__14843;
    wire N__14842;
    wire N__14839;
    wire N__14836;
    wire N__14833;
    wire N__14828;
    wire N__14825;
    wire N__14820;
    wire N__14819;
    wire N__14816;
    wire N__14813;
    wire N__14812;
    wire N__14807;
    wire N__14804;
    wire N__14799;
    wire N__14796;
    wire N__14793;
    wire N__14790;
    wire N__14787;
    wire N__14786;
    wire N__14785;
    wire N__14782;
    wire N__14777;
    wire N__14772;
    wire N__14771;
    wire N__14770;
    wire N__14767;
    wire N__14764;
    wire N__14759;
    wire N__14754;
    wire N__14753;
    wire N__14752;
    wire N__14749;
    wire N__14744;
    wire N__14739;
    wire N__14738;
    wire N__14737;
    wire N__14734;
    wire N__14731;
    wire N__14726;
    wire N__14721;
    wire N__14718;
    wire N__14715;
    wire N__14712;
    wire N__14709;
    wire N__14706;
    wire N__14703;
    wire N__14700;
    wire N__14697;
    wire N__14694;
    wire N__14693;
    wire N__14692;
    wire N__14691;
    wire N__14682;
    wire N__14679;
    wire N__14678;
    wire N__14675;
    wire N__14672;
    wire N__14671;
    wire N__14670;
    wire N__14661;
    wire N__14658;
    wire N__14655;
    wire N__14652;
    wire N__14651;
    wire N__14650;
    wire N__14647;
    wire N__14642;
    wire N__14637;
    wire N__14636;
    wire N__14635;
    wire N__14632;
    wire N__14629;
    wire N__14626;
    wire N__14623;
    wire N__14616;
    wire N__14615;
    wire N__14612;
    wire N__14611;
    wire N__14608;
    wire N__14603;
    wire N__14598;
    wire N__14597;
    wire N__14596;
    wire N__14593;
    wire N__14590;
    wire N__14587;
    wire N__14582;
    wire N__14577;
    wire N__14574;
    wire N__14571;
    wire N__14568;
    wire N__14565;
    wire N__14562;
    wire N__14559;
    wire N__14556;
    wire N__14553;
    wire N__14550;
    wire N__14547;
    wire N__14544;
    wire N__14541;
    wire N__14538;
    wire N__14535;
    wire N__14532;
    wire N__14529;
    wire N__14526;
    wire N__14525;
    wire N__14524;
    wire N__14521;
    wire N__14518;
    wire N__14515;
    wire N__14512;
    wire N__14509;
    wire N__14502;
    wire N__14501;
    wire N__14498;
    wire N__14497;
    wire N__14494;
    wire N__14491;
    wire N__14488;
    wire N__14481;
    wire N__14478;
    wire N__14475;
    wire N__14472;
    wire N__14469;
    wire N__14466;
    wire N__14463;
    wire N__14460;
    wire N__14457;
    wire N__14454;
    wire N__14451;
    wire N__14448;
    wire N__14445;
    wire N__14442;
    wire N__14439;
    wire GNDG0;
    wire VCCG0;
    wire CLK_c;
    wire \PWMInstance7.un1_periodCounter12_1_0_a2_0_6_cascade_ ;
    wire bfn_2_8_0_;
    wire \PWMInstance7.un1_periodCounter_2_cry_0 ;
    wire \PWMInstance7.un1_periodCounter_2_cry_1 ;
    wire \PWMInstance7.un1_periodCounter_2_cry_2 ;
    wire \PWMInstance7.un1_periodCounter_2_cry_3 ;
    wire \PWMInstance7.un1_periodCounter_2_cry_4 ;
    wire \PWMInstance7.un1_periodCounter_2_cry_5 ;
    wire \PWMInstance7.un1_periodCounter_2_cry_6 ;
    wire \PWMInstance7.un1_periodCounter_2_cry_7 ;
    wire bfn_2_9_0_;
    wire \PWMInstance7.un1_periodCounter_2_cry_8 ;
    wire \PWMInstance7.un1_periodCounter_2_cry_9 ;
    wire \PWMInstance7.un1_periodCounter_2_cry_10 ;
    wire \PWMInstance7.un1_periodCounter_2_cry_11 ;
    wire \PWMInstance7.un1_periodCounter_2_cry_12 ;
    wire \PWMInstance7.un1_periodCounter_2_cry_13 ;
    wire \PWMInstance7.un1_periodCounter_2_cry_14 ;
    wire \PWMInstance7.un1_periodCounter_2_cry_15 ;
    wire bfn_2_10_0_;
    wire \PWMInstance7.periodCounterZ0Z_16 ;
    wire \PWMInstance7.periodCounter12 ;
    wire \PWMInstance7.clkCountZ0Z_0 ;
    wire \PWMInstance7.clkCountZ0Z_1 ;
    wire \PWMInstance7.PWMPulseWidthCountZ0Z_2 ;
    wire \PWMInstance7.periodCounterZ0Z_2 ;
    wire \PWMInstance7.periodCounterZ0Z_3 ;
    wire \PWMInstance7.periodCounterZ0Z_11 ;
    wire \PWMInstance7.periodCounterZ0Z_10 ;
    wire \PWMInstance7.un1_periodCounter12_1_0_a2_0_0 ;
    wire \PWMInstance7.un1_periodCounter12_1_0_a2_0_10 ;
    wire \PWMInstance7.un1_periodCounter12_1_0_a2_0_9 ;
    wire \PWMInstance7.un1_periodCounter12_1_0_a2_0_12_cascade_ ;
    wire \PWMInstance7.un1_periodCounter12_1_0_a2_0_14 ;
    wire \PWMInstance7.periodCounterZ0Z_4 ;
    wire \PWMInstance7.periodCounterZ0Z_5 ;
    wire \PWMInstance7.periodCounterZ0Z_8 ;
    wire \PWMInstance7.periodCounterZ0Z_9 ;
    wire bfn_3_10_0_;
    wire \PWMInstance7.un1_PWMPulseWidthCount_0_I_9_c_RNO_6 ;
    wire \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_0 ;
    wire \PWMInstance7.un1_PWMPulseWidthCount_0_I_15_c_RNO_6 ;
    wire \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_1 ;
    wire \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_2 ;
    wire \PWMInstance7.un1_PWMPulseWidthCount_0_I_45_c_RNO_6 ;
    wire \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_3 ;
    wire \PWMInstance7.un1_PWMPulseWidthCount_0_I_33_c_RNO_6 ;
    wire \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_4 ;
    wire \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_5 ;
    wire \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_6 ;
    wire \PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_7 ;
    wire \PWMInstance7.un1_periodCounter12_1_0_a2_0 ;
    wire \PWMInstance7.out_0_sqmuxa ;
    wire bfn_3_11_0_;
    wire PWM7_c;
    wire pwmWrite_fastZ0Z_7;
    wire \PWMInstance7.PWMPulseWidthCountZ0Z_9 ;
    wire \PWMInstance7.PWMPulseWidthCountZ0Z_10 ;
    wire \PWMInstance7.PWMPulseWidthCountZ0Z_3 ;
    wire \PWMInstance7.periodCounterZ0Z_15 ;
    wire \PWMInstance7.periodCounterZ0Z_14 ;
    wire \PWMInstance7.un1_PWMPulseWidthCount_0_I_21_c_RNO_6 ;
    wire \PWMInstance7.PWMPulseWidthCountZ0Z_14 ;
    wire \PWMInstance7.periodCounterZ0Z_12 ;
    wire \PWMInstance7.periodCounterZ0Z_13 ;
    wire \PWMInstance7.un1_PWMPulseWidthCount_0_I_39_c_RNO_6 ;
    wire \PWMInstance7.periodCounterZ0Z_0 ;
    wire \PWMInstance7.periodCounterZ0Z_1 ;
    wire \PWMInstance7.un1_PWMPulseWidthCount_0_I_1_c_RNO_6 ;
    wire \PWMInstance7.periodCounterZ0Z_6 ;
    wire \PWMInstance7.periodCounterZ0Z_7 ;
    wire \PWMInstance7.un1_PWMPulseWidthCount_0_I_27_c_RNO_6 ;
    wire \PWMInstance7.PWMPulseWidthCountZ0Z_8 ;
    wire \PWMInstance7.PWMPulseWidthCountZ0Z_13 ;
    wire \PWMInstance7.PWMPulseWidthCountZ0Z_11 ;
    wire \PWMInstance7.PWMPulseWidthCountZ0Z_12 ;
    wire \PWMInstance7.PWMPulseWidthCountZ0Z_5 ;
    wire \PWMInstance7.PWMPulseWidthCountZ0Z_4 ;
    wire \PWMInstance7.PWMPulseWidthCountZ0Z_7 ;
    wire \PWMInstance7.PWMPulseWidthCountZ0Z_6 ;
    wire \PWMInstance7.PWMPulseWidthCountZ0Z_15 ;
    wire \PWMInstance7.PWMPulseWidthCountZ0Z_1 ;
    wire \PWMInstance7.PWMPulseWidthCountZ0Z_0 ;
    wire \PWMInstance7.pwmWrite_0_7 ;
    wire \PWMInstance5.PWMPulseWidthCountZ0Z_9 ;
    wire \PWMInstance5.PWMPulseWidthCountZ0Z_8 ;
    wire RST_c_i;
    wire ch0_B_c;
    wire \PWMInstance1.PWMPulseWidthCountZ0Z_2 ;
    wire \PWMInstance1.PWMPulseWidthCountZ0Z_3 ;
    wire \PWMInstance1.un1_periodCounter12_1_0_a2_0_0_cascade_ ;
    wire \PWMInstance1.PWMPulseWidthCountZ0Z_4 ;
    wire \PWMInstance1.PWMPulseWidthCountZ0Z_0 ;
    wire \PWMInstance1.PWMPulseWidthCountZ0Z_1 ;
    wire \PWMInstance1.PWMPulseWidthCountZ0Z_7 ;
    wire \PWMInstance1.PWMPulseWidthCountZ0Z_8 ;
    wire \PWMInstance1.PWMPulseWidthCountZ0Z_5 ;
    wire \PWMInstance1.PWMPulseWidthCountZ0Z_9 ;
    wire \PWMInstance1.PWMPulseWidthCountZ0Z_6 ;
    wire \PWMInstance1.PWMPulseWidthCountZ0Z_14 ;
    wire \PWMInstance1.PWMPulseWidthCountZ0Z_15 ;
    wire \PWMInstance1.PWMPulseWidthCountZ0Z_11 ;
    wire \PWMInstance1.PWMPulseWidthCountZ0Z_13 ;
    wire bfn_7_6_0_;
    wire \QuadInstance2.un1_Quad_cry_0 ;
    wire \QuadInstance2.un1_Quad_cry_1 ;
    wire \QuadInstance2.un1_Quad_cry_2 ;
    wire \QuadInstance2.un1_Quad_cry_3 ;
    wire \QuadInstance2.un1_Quad_cry_4 ;
    wire \QuadInstance2.un1_Quad_cry_5 ;
    wire \QuadInstance2.un1_Quad_cry_6 ;
    wire \QuadInstance2.un1_Quad_cry_7 ;
    wire bfn_7_7_0_;
    wire \QuadInstance2.un1_Quad_cry_8 ;
    wire \QuadInstance2.un1_Quad_cry_9 ;
    wire \QuadInstance2.un1_Quad_cry_10 ;
    wire \QuadInstance2.un1_Quad_cry_11 ;
    wire \QuadInstance2.un1_Quad_cry_12 ;
    wire \QuadInstance2.un1_Quad_cry_13 ;
    wire \QuadInstance2.un1_Quad_cry_14 ;
    wire \QuadInstance2.Quad_RNI8TLE2Z0Z_9 ;
    wire \QuadInstance2.Quad_RNIHU2G2Z0Z_11 ;
    wire \QuadInstance2.Quad_RNI0LLE2Z0Z_1 ;
    wire \QuadInstance2.Quad_RNIGT2G2Z0Z_10 ;
    wire \QuadInstance2.Quad_RNIIV2G2Z0Z_12 ;
    wire \QuadInstance2.Quad_RNI6RLE2Z0Z_7 ;
    wire \QuadInstance2.Quad_RNI7SLE2Z0Z_8 ;
    wire \QuadInstance2.Quad_RNI3OLE2Z0Z_4 ;
    wire \QuadInstance2.un1_Quad_axb_15 ;
    wire \QuadInstance2.count_enable_cascade_ ;
    wire \QuadInstance2.Quad_RNI1MLE2Z0Z_2 ;
    wire \QuadInstance2.un1_count_enable_i_a2_0_1_cascade_ ;
    wire \QuadInstance2.Quad_RNI2NLE2Z0Z_3 ;
    wire \QuadInstance2.Quad_RNI4PLE2Z0Z_5 ;
    wire \QuadInstance2.Quad_RNI5QLE2Z0Z_6 ;
    wire \QuadInstance2.delayedCh_AZ0Z_1 ;
    wire \QuadInstance2.delayedCh_AZ0Z_2 ;
    wire \QuadInstance2.Quad_RNIK13G2Z0Z_14 ;
    wire \QuadInstance2.delayedCh_BZ0Z_1 ;
    wire \QuadInstance2.delayedCh_BZ0Z_2 ;
    wire \PWMInstance1.un1_PWMPulseWidthCount_0_I_1_c_RNO_0 ;
    wire bfn_7_11_0_;
    wire \PWMInstance1.un1_PWMPulseWidthCount_0_I_9_c_RNO_0 ;
    wire \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_0 ;
    wire \PWMInstance1.un1_PWMPulseWidthCount_0_I_15_c_RNO_0 ;
    wire \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_1 ;
    wire \PWMInstance1.un1_PWMPulseWidthCount_0_I_27_c_RNO_0 ;
    wire \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_2 ;
    wire \PWMInstance1.un1_PWMPulseWidthCount_0_I_45_c_RNO_0 ;
    wire \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_3 ;
    wire \PWMInstance1.un1_PWMPulseWidthCount_0_I_33_c_RNO_0 ;
    wire \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_4 ;
    wire \PWMInstance1.un1_PWMPulseWidthCount_0_I_39_c_RNO_0 ;
    wire \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_5 ;
    wire \PWMInstance1.un1_PWMPulseWidthCount_0_I_21_c_RNO_0 ;
    wire \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_6 ;
    wire \PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_7 ;
    wire bfn_7_12_0_;
    wire PWM1_c;
    wire \PWMInstance0.PWMPulseWidthCountZ0Z_2 ;
    wire \PWMInstance0.PWMPulseWidthCountZ0Z_3 ;
    wire \PWMInstance0.un1_periodCounter12_1_0_a2_0_0_cascade_ ;
    wire \PWMInstance0.PWMPulseWidthCountZ0Z_5 ;
    wire \PWMInstance0.PWMPulseWidthCountZ0Z_4 ;
    wire pwmWrite_fastZ0Z_0;
    wire \PWMInstance0.clkCountZ0Z_1 ;
    wire \PWMInstance0.clkCountZ0Z_0 ;
    wire \PWMInstance0.periodCounter12_cascade_ ;
    wire \PWMInstance0.un1_periodCounter12_1_0_a2_0_6 ;
    wire \PWMInstance0.un1_periodCounter12_1_0_a2_0_10 ;
    wire \PWMInstance0.un1_periodCounter12_1_0_a2_0_14_cascade_ ;
    wire \PWMInstance0.un1_periodCounter12_1_0_a2_0_12 ;
    wire \PWMInstance0.periodCounter12 ;
    wire bfn_7_16_0_;
    wire \PWMInstance0.un1_periodCounter_2_cry_0 ;
    wire \PWMInstance0.periodCounterZ0Z_2 ;
    wire \PWMInstance0.un1_periodCounter_2_cry_1 ;
    wire \PWMInstance0.periodCounterZ0Z_3 ;
    wire \PWMInstance0.un1_periodCounter_2_cry_2 ;
    wire \PWMInstance0.periodCounterZ0Z_4 ;
    wire \PWMInstance0.un1_periodCounter_2_cry_3 ;
    wire \PWMInstance0.periodCounterZ0Z_5 ;
    wire \PWMInstance0.un1_periodCounter_2_cry_4 ;
    wire \PWMInstance0.un1_periodCounter_2_cry_5 ;
    wire \PWMInstance0.un1_periodCounter_2_cry_6 ;
    wire \PWMInstance0.un1_periodCounter_2_cry_7 ;
    wire bfn_7_17_0_;
    wire \PWMInstance0.un1_periodCounter_2_cry_8 ;
    wire \PWMInstance0.un1_periodCounter_2_cry_9 ;
    wire \PWMInstance0.un1_periodCounter_2_cry_10 ;
    wire \PWMInstance0.un1_periodCounter_2_cry_11 ;
    wire \PWMInstance0.un1_periodCounter_2_cry_12 ;
    wire \PWMInstance0.un1_periodCounter_2_cry_13 ;
    wire \PWMInstance0.un1_periodCounter_2_cry_14 ;
    wire \PWMInstance0.un1_periodCounter_2_cry_15 ;
    wire bfn_7_18_0_;
    wire \PWMInstance0.periodCounterZ0Z_16 ;
    wire \PWMInstance1.periodCounterZ0Z_0 ;
    wire bfn_8_1_0_;
    wire \PWMInstance1.un1_periodCounter_2_cry_0 ;
    wire \PWMInstance1.periodCounterZ0Z_2 ;
    wire \PWMInstance1.un1_periodCounter_2_cry_1 ;
    wire \PWMInstance1.periodCounterZ0Z_3 ;
    wire \PWMInstance1.un1_periodCounter_2_cry_2 ;
    wire \PWMInstance1.periodCounterZ0Z_4 ;
    wire \PWMInstance1.un1_periodCounter_2_cry_3 ;
    wire \PWMInstance1.periodCounterZ0Z_5 ;
    wire \PWMInstance1.un1_periodCounter_2_cry_4 ;
    wire \PWMInstance1.periodCounterZ0Z_6 ;
    wire \PWMInstance1.un1_periodCounter_2_cry_5 ;
    wire \PWMInstance1.un1_periodCounter_2_cry_6 ;
    wire \PWMInstance1.un1_periodCounter_2_cry_7 ;
    wire \PWMInstance1.periodCounterZ0Z_8 ;
    wire bfn_8_2_0_;
    wire \PWMInstance1.periodCounterZ0Z_9 ;
    wire \PWMInstance1.un1_periodCounter_2_cry_8 ;
    wire \PWMInstance1.periodCounterZ0Z_10 ;
    wire \PWMInstance1.un1_periodCounter_2_cry_9 ;
    wire \PWMInstance1.periodCounterZ0Z_11 ;
    wire \PWMInstance1.un1_periodCounter_2_cry_10 ;
    wire \PWMInstance1.periodCounterZ0Z_12 ;
    wire \PWMInstance1.un1_periodCounter_2_cry_11 ;
    wire \PWMInstance1.periodCounterZ0Z_13 ;
    wire \PWMInstance1.un1_periodCounter_2_cry_12 ;
    wire \PWMInstance1.periodCounterZ0Z_14 ;
    wire \PWMInstance1.un1_periodCounter_2_cry_13 ;
    wire \PWMInstance1.un1_periodCounter_2_cry_14 ;
    wire \PWMInstance1.un1_periodCounter_2_cry_15 ;
    wire bfn_8_3_0_;
    wire bfn_8_4_0_;
    wire \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_0 ;
    wire \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_1 ;
    wire \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_2 ;
    wire \PWMInstance5.un1_PWMPulseWidthCount_0_I_45_c_RNO_4 ;
    wire \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_3 ;
    wire \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_4 ;
    wire \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_5 ;
    wire \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_6 ;
    wire \PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_7 ;
    wire bfn_8_5_0_;
    wire PWM5_c;
    wire \PWMInstance1.PWMPulseWidthCountZ0Z_12 ;
    wire \PWMInstance1.PWMPulseWidthCountZ0Z_10 ;
    wire \QuadInstance2.Quad_RNO_0_2_9 ;
    wire \QuadInstance2.Quad_RNO_0_2_10 ;
    wire \QuadInstance2.Quad_RNO_0_2_14 ;
    wire \QuadInstance2.Quad_RNO_0_2_12 ;
    wire \QuadInstance7.un1_count_enable_i_a2_0_1_cascade_ ;
    wire \QuadInstance7.count_enable_cascade_ ;
    wire \QuadInstance7.un1_count_enable_i_a2_0_1 ;
    wire \QuadInstance7.delayedCh_AZ0Z_1 ;
    wire \QuadInstance7.delayedCh_AZ0Z_2 ;
    wire \QuadInstance7.delayedCh_BZ0Z_1 ;
    wire \QuadInstance7.delayedCh_BZ0Z_2 ;
    wire \PWMInstance1.un1_periodCounter12_1_0_a2_0 ;
    wire \PWMInstance1.pwmWrite_0_1 ;
    wire pwmWriteZ0Z_1;
    wire \PWMInstance1.clkCountZ0Z_1 ;
    wire \PWMInstance1.clkCountZ0Z_0 ;
    wire \PWMInstance1.periodCounterZ0Z_16 ;
    wire \PWMInstance1.periodCounterZ0Z_7 ;
    wire \PWMInstance1.periodCounterZ0Z_15 ;
    wire \PWMInstance1.periodCounterZ0Z_1 ;
    wire \PWMInstance1.un1_periodCounter12_1_0_a2_0_6_cascade_ ;
    wire \PWMInstance1.periodCounter12 ;
    wire \PWMInstance1.un1_periodCounter12_1_0_a2_0_10 ;
    wire \PWMInstance1.un1_periodCounter12_1_0_a2_0_9 ;
    wire \PWMInstance1.un1_periodCounter12_1_0_a2_0_14_cascade_ ;
    wire \PWMInstance1.un1_periodCounter12_1_0_a2_0_12 ;
    wire \PWMInstance1.out_0_sqmuxa ;
    wire \PWMInstance5.un1_PWMPulseWidthCount_0_I_9_c_RNO_4 ;
    wire \PWMInstance5.PWMPulseWidthCountZ0Z_2 ;
    wire \PWMInstance5.PWMPulseWidthCountZ0Z_3 ;
    wire \PWMInstance5.PWMPulseWidthCountZ0Z_14 ;
    wire \PWMInstance5.un1_PWMPulseWidthCount_0_I_21_c_RNO_4 ;
    wire \PWMInstance5.PWMPulseWidthCountZ0Z_15 ;
    wire \PWMInstance0.PWMPulseWidthCountZ0Z_9 ;
    wire \PWMInstance0.periodCounterZ0Z_9 ;
    wire \PWMInstance0.PWMPulseWidthCountZ0Z_8 ;
    wire pwmWriteZ0Z_0;
    wire \PWMInstance5.PWMPulseWidthCountZ0Z_12 ;
    wire \PWMInstance5.un1_PWMPulseWidthCount_0_I_39_c_RNO_4 ;
    wire \PWMInstance0.PWMPulseWidthCountZ0Z_6 ;
    wire \PWMInstance0.periodCounterZ0Z_7 ;
    wire \PWMInstance0.periodCounterZ0Z_15 ;
    wire \PWMInstance0.periodCounterZ0Z_14 ;
    wire \PWMInstance0.PWMPulseWidthCountZ0Z_14 ;
    wire \PWMInstance0.PWMPulseWidthCountZ0Z_15 ;
    wire \PWMInstance0.periodCounterZ0Z_10 ;
    wire \PWMInstance0.periodCounterZ0Z_11 ;
    wire \PWMInstance0.PWMPulseWidthCountZ0Z_10 ;
    wire \PWMInstance0.PWMPulseWidthCountZ0Z_11 ;
    wire \PWMInstance0.PWMPulseWidthCountZ0Z_13 ;
    wire \PWMInstance0.PWMPulseWidthCountZ0Z_12 ;
    wire \PWMInstance0.periodCounterZ0Z_12 ;
    wire bfn_8_15_0_;
    wire \PWMInstance0.un1_PWMPulseWidthCount_0_I_9_c_RNOZ0 ;
    wire \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_0 ;
    wire \PWMInstance0.un1_PWMPulseWidthCount_0_I_15_c_RNOZ0 ;
    wire \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_1 ;
    wire \PWMInstance0.un1_PWMPulseWidthCount_0_I_27_c_RNOZ0 ;
    wire \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_2 ;
    wire \PWMInstance0.un1_PWMPulseWidthCount_0_I_45_c_RNOZ0 ;
    wire \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_3 ;
    wire \PWMInstance0.un1_PWMPulseWidthCount_0_I_33_c_RNOZ0 ;
    wire \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_4 ;
    wire \PWMInstance0.un1_PWMPulseWidthCount_0_I_39_c_RNOZ0 ;
    wire \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_5 ;
    wire \PWMInstance0.un1_PWMPulseWidthCount_0_I_21_c_RNOZ0 ;
    wire \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_6 ;
    wire \PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_7 ;
    wire \PWMInstance0.un1_periodCounter12_1_0_a2_0 ;
    wire \PWMInstance0.out_0_sqmuxa ;
    wire bfn_8_16_0_;
    wire PWM0_c;
    wire ch7_B_c;
    wire \QuadInstance7.delayedCh_BZ0Z_0 ;
    wire PWM0_obufLegalizeSB_DFFNet;
    wire PWM1_obufLegalizeSB_DFFNet;
    wire PWM6_obufLegalizeSB_DFFNet;
    wire PWM7_obufLegalizeSB_DFFNet;
    wire ch3_B_c;
    wire \QuadInstance2.Quad_RNO_0_2_4 ;
    wire ch5_A_c;
    wire \QuadInstance5.delayedCh_AZ0Z_0 ;
    wire \QuadInstance5.un1_count_enable_i_a2_0_1_cascade_ ;
    wire \QuadInstance2.un1_count_enable_i_a2_0_1 ;
    wire \QuadInstance2.Quad_RNIJ03G2Z0Z_13 ;
    wire \QuadInstance5.un1_count_enable_i_a2_0_1 ;
    wire bfn_9_8_0_;
    wire \QuadInstance7.Quad_RNI85VV2Z0Z_1 ;
    wire \QuadInstance7.un1_Quad_cry_0 ;
    wire \QuadInstance7.Quad_RNI96VV2Z0Z_2 ;
    wire \QuadInstance7.un1_Quad_cry_1 ;
    wire \QuadInstance7.Quad_RNIA7VV2Z0Z_3 ;
    wire \QuadInstance7.un1_Quad_cry_2 ;
    wire \QuadInstance7.Quad_RNIB8VV2Z0Z_4 ;
    wire \QuadInstance7.un1_Quad_cry_3 ;
    wire \QuadInstance7.Quad_RNIC9VV2Z0Z_5 ;
    wire \QuadInstance7.un1_Quad_cry_4 ;
    wire \QuadInstance7.Quad_RNIDAVV2Z0Z_6 ;
    wire \QuadInstance7.un1_Quad_cry_5 ;
    wire \QuadInstance7.Quad_RNIEBVV2Z0Z_7 ;
    wire \QuadInstance7.un1_Quad_cry_6 ;
    wire \QuadInstance7.un1_Quad_cry_7 ;
    wire \QuadInstance7.Quad_RNIFCVV2Z0Z_8 ;
    wire bfn_9_9_0_;
    wire \QuadInstance7.Quad_RNIGDVV2Z0Z_9 ;
    wire \QuadInstance7.un1_Quad_cry_8 ;
    wire \QuadInstance7.Quad_RNIOIKU2Z0Z_10 ;
    wire \QuadInstance7.un1_Quad_cry_9 ;
    wire \QuadInstance7.Quad_RNIPJKU2Z0Z_11 ;
    wire \QuadInstance7.Quad_RNO_0_7_11 ;
    wire \QuadInstance7.un1_Quad_cry_10 ;
    wire \QuadInstance7.Quad_RNIQKKU2Z0Z_12 ;
    wire \QuadInstance7.Quad_RNO_0_7_12 ;
    wire \QuadInstance7.un1_Quad_cry_11 ;
    wire \QuadInstance7.Quad_RNIRLKU2Z0Z_13 ;
    wire \QuadInstance7.un1_Quad_cry_12 ;
    wire \QuadInstance7.Quad_RNISMKU2Z0Z_14 ;
    wire \QuadInstance7.un1_Quad_cry_13 ;
    wire \QuadInstance7.un1_Quad_axb_15 ;
    wire \QuadInstance7.un1_Quad_cry_14 ;
    wire pwmWrite_fastZ0Z_1;
    wire pwmWriteZ0Z_7;
    wire \PWMInstance5.un1_PWMPulseWidthCount_0_I_1_c_RNO_4 ;
    wire \PWMInstance5.PWMPulseWidthCountZ0Z_0 ;
    wire \PWMInstance5.PWMPulseWidthCountZ0Z_1 ;
    wire \PWMInstance5.un1_PWMPulseWidthCount_0_I_27_c_RNO_4 ;
    wire \PWMInstance5.PWMPulseWidthCountZ0Z_6 ;
    wire \PWMInstance5.PWMPulseWidthCountZ0Z_7 ;
    wire \PWMInstance5.periodCounterZ0Z_0 ;
    wire bfn_9_12_0_;
    wire \PWMInstance5.un1_periodCounter_2_cry_0 ;
    wire \PWMInstance5.un1_periodCounter_2_cry_1 ;
    wire \PWMInstance5.un1_periodCounter_2_cry_2 ;
    wire \PWMInstance5.un1_periodCounter_2_cry_3 ;
    wire \PWMInstance5.un1_periodCounter_2_cry_4 ;
    wire \PWMInstance5.periodCounterZ0Z_6 ;
    wire \PWMInstance5.un1_periodCounter_2_cry_5 ;
    wire \PWMInstance5.un1_periodCounter_2_cry_6 ;
    wire \PWMInstance5.un1_periodCounter_2_cry_7 ;
    wire \PWMInstance5.periodCounterZ0Z_8 ;
    wire bfn_9_13_0_;
    wire \PWMInstance5.un1_periodCounter_2_cry_8 ;
    wire \PWMInstance5.un1_periodCounter_2_cry_9 ;
    wire \PWMInstance5.un1_periodCounter_2_cry_10 ;
    wire \PWMInstance5.un1_periodCounter_2_cry_11 ;
    wire \PWMInstance5.periodCounterZ0Z_13 ;
    wire \PWMInstance5.un1_periodCounter_2_cry_12 ;
    wire \PWMInstance5.un1_periodCounter_2_cry_13 ;
    wire \PWMInstance5.un1_periodCounter_2_cry_14 ;
    wire \PWMInstance5.un1_periodCounter_2_cry_15 ;
    wire bfn_9_14_0_;
    wire \PWMInstance0.periodCounterZ0Z_8 ;
    wire \PWMInstance0.periodCounterZ0Z_6 ;
    wire \PWMInstance0.periodCounterZ0Z_13 ;
    wire \PWMInstance0.un1_periodCounter12_1_0_a2_0_9 ;
    wire \PWMInstance0.periodCounterZ0Z_0 ;
    wire \PWMInstance0.periodCounterZ0Z_1 ;
    wire \PWMInstance0.un1_PWMPulseWidthCount_0_I_1_c_RNOZ0 ;
    wire \PWMInstance0.PWMPulseWidthCountZ0Z_0 ;
    wire \PWMInstance0.PWMPulseWidthCountZ0Z_1 ;
    wire \PWMInstance0.PWMPulseWidthCountZ0Z_7 ;
    wire \PWMInstance0.pwmWrite_0_0 ;
    wire \PWMInstance5.PWMPulseWidthCountZ0Z_13 ;
    wire ch5_B_c;
    wire \QuadInstance5.delayedCh_BZ0Z_0 ;
    wire \QuadInstance2.count_enable ;
    wire \QuadInstance5.delayedCh_BZ0Z_1 ;
    wire \QuadInstance5.delayedCh_AZ0Z_1 ;
    wire \QuadInstance5.delayedCh_AZ0Z_2 ;
    wire \QuadInstance5.delayedCh_BZ0Z_2 ;
    wire \QuadInstance5.count_enable_cascade_ ;
    wire \QuadInstance5.count_enable ;
    wire bfn_10_6_0_;
    wire \QuadInstance5.Quad_RNIOUKI2Z0Z_1 ;
    wire \QuadInstance5.Quad_RNO_0_4_1 ;
    wire \QuadInstance5.un1_Quad_cry_0 ;
    wire \QuadInstance5.Quad_RNIPVKI2Z0Z_2 ;
    wire \QuadInstance5.un1_Quad_cry_1 ;
    wire \QuadInstance5.Quad_RNIQ0LI2Z0Z_3 ;
    wire \QuadInstance5.un1_Quad_cry_2 ;
    wire \QuadInstance5.Quad_RNIR1LI2Z0Z_4 ;
    wire \QuadInstance5.un1_Quad_cry_3 ;
    wire \QuadInstance5.Quad_RNIS2LI2Z0Z_5 ;
    wire \QuadInstance5.un1_Quad_cry_4 ;
    wire \QuadInstance5.Quad_RNIT3LI2Z0Z_6 ;
    wire \QuadInstance5.un1_Quad_cry_5 ;
    wire \QuadInstance5.Quad_RNIU4LI2Z0Z_7 ;
    wire \QuadInstance5.un1_Quad_cry_6 ;
    wire \QuadInstance5.un1_Quad_cry_7 ;
    wire \QuadInstance5.Quad_RNIV5LI2Z0Z_8 ;
    wire bfn_10_7_0_;
    wire \QuadInstance5.Quad_RNI07LI2Z0Z_9 ;
    wire \QuadInstance5.un1_Quad_cry_8 ;
    wire \QuadInstance5.Quad_RNI8AQ82Z0Z_10 ;
    wire \QuadInstance5.un1_Quad_cry_9 ;
    wire \QuadInstance5.Quad_RNI9BQ82Z0Z_11 ;
    wire \QuadInstance5.un1_Quad_cry_10 ;
    wire \QuadInstance5.Quad_RNIACQ82Z0Z_12 ;
    wire \QuadInstance5.Quad_RNO_0_5_12 ;
    wire \QuadInstance5.un1_Quad_cry_11 ;
    wire \QuadInstance5.Quad_RNIBDQ82Z0Z_13 ;
    wire \QuadInstance5.Quad_RNO_0_5_13 ;
    wire \QuadInstance5.un1_Quad_cry_12 ;
    wire \QuadInstance5.Quad_RNICEQ82Z0Z_14 ;
    wire \QuadInstance5.Quad_RNO_0_5_14 ;
    wire \QuadInstance5.un1_Quad_cry_13 ;
    wire \QuadInstance5.un1_Quad_axb_15 ;
    wire \QuadInstance5.un1_Quad_cry_14 ;
    wire bfn_10_8_0_;
    wire \QuadInstance3.un1_Quad_cry_0 ;
    wire \QuadInstance3.un1_Quad_cry_1 ;
    wire \QuadInstance3.Quad_RNIAQAL1Z0Z_3 ;
    wire \QuadInstance3.un1_Quad_cry_2 ;
    wire \QuadInstance3.un1_Quad_cry_3 ;
    wire \QuadInstance3.Quad_RNICSAL1Z0Z_5 ;
    wire \QuadInstance3.un1_Quad_cry_4 ;
    wire \QuadInstance3.Quad_RNIDTAL1Z0Z_6 ;
    wire \QuadInstance3.un1_Quad_cry_5 ;
    wire \QuadInstance3.un1_Quad_cry_6 ;
    wire \QuadInstance3.un1_Quad_cry_7 ;
    wire bfn_10_9_0_;
    wire \QuadInstance3.un1_Quad_cry_8 ;
    wire \QuadInstance3.un1_Quad_cry_9 ;
    wire \QuadInstance3.Quad_RNIP20J1Z0Z_11 ;
    wire \QuadInstance3.un1_Quad_cry_10 ;
    wire \QuadInstance3.Quad_RNIQ30J1Z0Z_12 ;
    wire \QuadInstance3.un1_Quad_cry_11 ;
    wire \QuadInstance3.Quad_RNIR40J1Z0Z_13 ;
    wire \QuadInstance3.un1_Quad_cry_12 ;
    wire \QuadInstance3.un1_Quad_cry_13 ;
    wire \QuadInstance3.un1_Quad_cry_14 ;
    wire \QuadInstance3.count_enable_cascade_ ;
    wire \QuadInstance3.Quad_RNI8OAL1Z0Z_1 ;
    wire \QuadInstance3.un1_count_enable_i_a2_0_1_cascade_ ;
    wire \QuadInstance3.Quad_RNI9PAL1Z0Z_2 ;
    wire \QuadInstance3.Quad_RNIO10J1Z0Z_10 ;
    wire \QuadInstance3.Quad_RNIFVAL1Z0Z_8 ;
    wire \QuadInstance3.Quad_RNIG0BL1Z0Z_9 ;
    wire \QuadInstance3.Quad_RNIBRAL1Z0Z_4 ;
    wire \QuadInstance3.Quad_RNIS50J1Z0Z_14 ;
    wire \QuadInstance3.delayedCh_BZ0Z_2 ;
    wire \QuadInstance3.delayedCh_AZ0Z_2 ;
    wire \QuadInstance3.delayedCh_AZ0Z_1 ;
    wire \QuadInstance3.Quad_RNIEUAL1Z0Z_7 ;
    wire \QuadInstance3.un1_count_enable_i_a2_0_1 ;
    wire \QuadInstance3.count_enable ;
    wire \QuadInstance3.un1_Quad_axb_15 ;
    wire \QuadInstance3.delayedCh_BZ0Z_0 ;
    wire \QuadInstance3.delayedCh_BZ0Z_1 ;
    wire \PWMInstance5.un1_PWMPulseWidthCount_0_I_15_c_RNO_4 ;
    wire \PWMInstance5.periodCounterZ0Z_2 ;
    wire \PWMInstance5.periodCounterZ0Z_14 ;
    wire \PWMInstance5.periodCounterZ0Z_12 ;
    wire \PWMInstance5.un1_periodCounter12_1_0_a2_0_0_cascade_ ;
    wire \PWMInstance5.periodCounterZ0Z_4 ;
    wire \PWMInstance5.PWMPulseWidthCountZ0Z_4 ;
    wire \PWMInstance5.PWMPulseWidthCountZ0Z_5 ;
    wire \PWMInstance5.periodCounterZ0Z_10 ;
    wire \PWMInstance5.PWMPulseWidthCountZ0Z_10 ;
    wire \PWMInstance5.un1_PWMPulseWidthCount_0_I_33_c_RNO_4 ;
    wire \PWMInstance5.PWMPulseWidthCountZ0Z_11 ;
    wire \PWMInstance5.un1_periodCounter12_1_0_a2_0 ;
    wire \PWMInstance5.pwmWrite_0_5 ;
    wire \PWMInstance5.clkCountZ0Z_1 ;
    wire \PWMInstance5.clkCountZ0Z_0 ;
    wire \PWMInstance5.periodCounter12 ;
    wire \PWMInstance5.periodCounterZ0Z_15 ;
    wire \PWMInstance5.periodCounterZ0Z_1 ;
    wire \PWMInstance5.periodCounter12_cascade_ ;
    wire \PWMInstance5.un1_periodCounter12_1_0_a2_0_9 ;
    wire \PWMInstance5.un1_periodCounter12_1_0_a2_0_14_cascade_ ;
    wire \PWMInstance5.un1_periodCounter12_1_0_a2_0_12 ;
    wire \PWMInstance5.out_0_sqmuxa ;
    wire \PWMInstance5.periodCounterZ0Z_9 ;
    wire \PWMInstance5.periodCounterZ0Z_5 ;
    wire \PWMInstance5.periodCounterZ0Z_11 ;
    wire \PWMInstance5.periodCounterZ0Z_3 ;
    wire \PWMInstance5.un1_periodCounter12_1_0_a2_0_10 ;
    wire \PWMInstance5.periodCounterZ0Z_16 ;
    wire \PWMInstance5.periodCounterZ0Z_7 ;
    wire \PWMInstance5.un1_periodCounter12_1_0_a2_0_6 ;
    wire \PWMInstance6.un1_periodCounter12_1_0_a2_0_0_cascade_ ;
    wire \PWMInstance6.un1_periodCounter12_1_0_a2_0_12_cascade_ ;
    wire \PWMInstance6.un1_periodCounter12_1_0_a2_0_10 ;
    wire \PWMInstance6.PWMPulseWidthCountZ0Z_2 ;
    wire \PWMInstance6.PWMPulseWidthCountZ0Z_3 ;
    wire \PWMInstance6.PWMPulseWidthCountZ0Z_4 ;
    wire \QuadInstance2.Quad_RNO_0_2_2 ;
    wire \QuadInstance3.Quad_RNO_0_3_2 ;
    wire \QuadInstance2.Quad_RNO_0_2_6 ;
    wire \QuadInstance7.Quad_RNO_0_7_2 ;
    wire \QuadInstance2.Quad_RNO_0_2_3 ;
    wire \QuadInstance5.Quad_RNO_0_5_4 ;
    wire \QuadInstance5.Quad_RNO_0_5_6 ;
    wire \QuadInstance7.Quad_RNO_0_7_6 ;
    wire \QuadInstance7.Quad_RNO_0_7_9 ;
    wire \QuadInstance5.Quad_RNO_0_5_8 ;
    wire \QuadInstance3.Quad_RNO_0_3_3 ;
    wire \QuadInstance2.Quad_RNO_0_2_7 ;
    wire \QuadInstance3.Quad_RNO_0_3_7 ;
    wire \QuadInstance5.Quad_RNO_0_5_7 ;
    wire \QuadInstance3.Quad_RNO_0_3_5 ;
    wire \QuadInstance7.Quad_RNO_0_7_7 ;
    wire \QuadInstance2.Quad_RNO_0_2_11 ;
    wire \QuadInstance5.Quad_RNO_0_5_10 ;
    wire \QuadInstance5.Quad_RNO_0_5_11 ;
    wire \QuadInstance2.Quad_RNO_0_2_8 ;
    wire \QuadInstance3.Quad_RNO_0_3_9 ;
    wire dataRead5_13;
    wire \QuadInstance2.Quad_RNO_0_2_13 ;
    wire dataRead2_13;
    wire \QuadInstance3.Quad_RNO_0_3_13 ;
    wire dataRead3_13;
    wire \QuadInstance3.Quad_RNO_0_3_12 ;
    wire \QuadInstance3.Quad_RNO_0_3_8 ;
    wire \QuadInstance3.Quad_RNO_0_3_14 ;
    wire \QuadInstance5.Quad_RNO_0_5_2 ;
    wire \QuadInstance7.Quad_RNO_0_7_14 ;
    wire \QuadInstance3.Quad_RNO_0_3_10 ;
    wire \QuadInstance3.Quad_RNO_0_3_11 ;
    wire OutReg_ess_RNO_2Z0Z_13;
    wire dataRead5_11;
    wire OutReg_0_5_i_m3_i_m3_ns_1_11_cascade_;
    wire dataRead3_14;
    wire dataRead2_14;
    wire dataRead7_14;
    wire OutReg_0_4_i_m3_ns_1_14_cascade_;
    wire pwmWrite_fastZ0Z_5;
    wire pwmWriteZ0Z_5;
    wire bfn_11_14_0_;
    wire \PWMInstance6.un1_periodCounter_2_cry_0 ;
    wire \PWMInstance6.periodCounterZ0Z_2 ;
    wire \PWMInstance6.un1_periodCounter_2_cry_1 ;
    wire \PWMInstance6.periodCounterZ0Z_3 ;
    wire \PWMInstance6.un1_periodCounter_2_cry_2 ;
    wire \PWMInstance6.periodCounterZ0Z_4 ;
    wire \PWMInstance6.un1_periodCounter_2_cry_3 ;
    wire \PWMInstance6.periodCounterZ0Z_5 ;
    wire \PWMInstance6.un1_periodCounter_2_cry_4 ;
    wire \PWMInstance6.un1_periodCounter_2_cry_5 ;
    wire \PWMInstance6.un1_periodCounter_2_cry_6 ;
    wire \PWMInstance6.un1_periodCounter_2_cry_7 ;
    wire bfn_11_15_0_;
    wire \PWMInstance6.un1_periodCounter_2_cry_8 ;
    wire \PWMInstance6.un1_periodCounter_2_cry_9 ;
    wire \PWMInstance6.un1_periodCounter_2_cry_10 ;
    wire \PWMInstance6.un1_periodCounter_2_cry_11 ;
    wire \PWMInstance6.un1_periodCounter_2_cry_12 ;
    wire \PWMInstance6.un1_periodCounter_2_cry_13 ;
    wire \PWMInstance6.un1_periodCounter_2_cry_14 ;
    wire \PWMInstance6.un1_periodCounter_2_cry_15 ;
    wire bfn_11_16_0_;
    wire ch3_A_c;
    wire \QuadInstance3.delayedCh_AZ0Z_0 ;
    wire \QuadInstance2.Quad_RNO_0_2_5 ;
    wire \QuadInstance5.Quad_RNO_0_5_5 ;
    wire \QuadInstance7.Quad_RNO_0_7_5 ;
    wire bfn_12_5_0_;
    wire \QuadInstance6.un1_Quad_cry_0 ;
    wire \QuadInstance6.Quad_RNO_0_6_2 ;
    wire \QuadInstance6.un1_Quad_cry_1 ;
    wire \QuadInstance6.Quad_RNO_0_6_3 ;
    wire \QuadInstance6.un1_Quad_cry_2 ;
    wire \QuadInstance6.un1_Quad_cry_3 ;
    wire \QuadInstance6.Quad_RNO_0_6_5 ;
    wire \QuadInstance6.un1_Quad_cry_4 ;
    wire \QuadInstance6.Quad_RNO_0_6_6 ;
    wire \QuadInstance6.un1_Quad_cry_5 ;
    wire \QuadInstance6.Quad_RNO_0_6_7 ;
    wire \QuadInstance6.un1_Quad_cry_6 ;
    wire \QuadInstance6.un1_Quad_cry_7 ;
    wire \QuadInstance6.Quad_RNO_0_6_8 ;
    wire bfn_12_6_0_;
    wire \QuadInstance6.un1_Quad_cry_8 ;
    wire \QuadInstance6.un1_Quad_cry_9 ;
    wire \QuadInstance6.Quad_RNO_0_6_11 ;
    wire \QuadInstance6.un1_Quad_cry_10 ;
    wire \QuadInstance6.Quad_RNO_0_6_12 ;
    wire \QuadInstance6.un1_Quad_cry_11 ;
    wire \QuadInstance6.Quad_RNO_0_6_13 ;
    wire \QuadInstance6.un1_Quad_cry_12 ;
    wire \QuadInstance6.Quad_RNIKINB1Z0Z_14 ;
    wire \QuadInstance6.un1_Quad_cry_13 ;
    wire \QuadInstance6.un1_Quad_axb_15 ;
    wire \QuadInstance6.un1_Quad_cry_14 ;
    wire \QuadInstance6.Quad_RNO_0_5_1 ;
    wire \QuadInstance7.Quad_RNO_0_7_8 ;
    wire \QuadInstance6.Quad_RNO_0_6_14 ;
    wire dataRead6_14;
    wire \QuadInstance6.Quad_RNO_0_6_10 ;
    wire \QuadInstance7.Quad_RNO_0_7_10 ;
    wire \QuadInstance5.Quad_RNO_0_5_9 ;
    wire \QuadInstance6.Quad_RNI02A91Z0Z_1 ;
    wire \QuadInstance6.count_enable_cascade_ ;
    wire \QuadInstance6.Quad_RNI13A91Z0Z_2 ;
    wire \QuadInstance6.Quad_RNIHFNB1Z0Z_11 ;
    wire \QuadInstance6.Quad_RNI24A91Z0Z_3 ;
    wire \QuadInstance6.Quad_RNI46A91Z0Z_5 ;
    wire \QuadInstance6.Quad_RNI8AA91Z0Z_9 ;
    wire \QuadInstance6.Quad_RNI79A91Z0Z_8 ;
    wire \QuadInstance6.un1_count_enable_i_a2_0_1_cascade_ ;
    wire \QuadInstance6.Quad_RNI35A91Z0Z_4 ;
    wire \QuadInstance6.Quad_RNIIGNB1Z0Z_12 ;
    wire \QuadInstance6.Quad_RNI57A91Z0Z_6 ;
    wire \QuadInstance6.Quad_RNI68A91Z0Z_7 ;
    wire OutReg_0_4_i_m3_ns_1_13;
    wire OutReg_ess_RNO_1Z0Z_13;
    wire dataRead7_11;
    wire dataRead6_11;
    wire OutReg_ess_RNO_1Z0Z_11_cascade_;
    wire OutReg_ess_RNO_2Z0Z_11;
    wire OutReg_ess_RNO_0Z0Z_11_cascade_;
    wire OutReg_ess_RNO_0Z0Z_13;
    wire data_receivedZ0Z_18;
    wire data_receivedZ0Z_17;
    wire data_receivedZ0Z_16;
    wire data_receivedZ0Z_15;
    wire \PWMInstance6.clkCountZ0Z_0 ;
    wire \PWMInstance6.clkCountZ0Z_1 ;
    wire pwmWrite_fastZ0Z_6;
    wire pwmWriteZ0Z_6;
    wire \PWMInstance6.periodCounterZ0Z_16 ;
    wire \PWMInstance6.un1_periodCounter12_1_0_a2_0_6_cascade_ ;
    wire \PWMInstance6.periodCounter12 ;
    wire \PWMInstance6.un1_periodCounter12_1_0_a2_0_14 ;
    wire ch6_A_c;
    wire \QuadInstance6.delayedCh_AZ0Z_0 ;
    wire \PWMInstance6.un1_periodCounter12_1_0_a2_0_9 ;
    wire \PWMInstance6.periodCounterZ0Z_0 ;
    wire \PWMInstance6.periodCounterZ0Z_1 ;
    wire \PWMInstance6.PWMPulseWidthCountZ0Z_0 ;
    wire \PWMInstance6.PWMPulseWidthCountZ0Z_1 ;
    wire \PWMInstance6.periodCounterZ0Z_6 ;
    wire \PWMInstance6.periodCounterZ0Z_7 ;
    wire \PWMInstance6.PWMPulseWidthCountZ0Z_6 ;
    wire \PWMInstance6.PWMPulseWidthCountZ0Z_7 ;
    wire \PWMInstance6.periodCounterZ0Z_8 ;
    wire \PWMInstance6.periodCounterZ0Z_9 ;
    wire \PWMInstance6.un1_PWMPulseWidthCount_0_I_1_c_RNO_5 ;
    wire bfn_12_16_0_;
    wire \PWMInstance6.un1_PWMPulseWidthCount_0_I_9_c_RNO_5 ;
    wire \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_0 ;
    wire \PWMInstance6.un1_PWMPulseWidthCount_0_I_15_c_RNO_5 ;
    wire \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_1 ;
    wire \PWMInstance6.un1_PWMPulseWidthCount_0_I_27_c_RNO_5 ;
    wire \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_2 ;
    wire \PWMInstance6.un1_PWMPulseWidthCount_0_I_45_c_RNO_5 ;
    wire \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_3 ;
    wire \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_4 ;
    wire \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_5 ;
    wire \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_6 ;
    wire \PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_7 ;
    wire \PWMInstance6.un1_periodCounter12_1_0_a2_0 ;
    wire \PWMInstance6.out_0_sqmuxa ;
    wire bfn_12_17_0_;
    wire PWM6_c;
    wire PWM5_obufLegalizeSB_DFFNet;
    wire ch2_A_c;
    wire \QuadInstance2.delayedCh_AZ0Z_0 ;
    wire dataRead5_4;
    wire OutReg_ess_RNO_2Z0Z_4_cascade_;
    wire dataRead2_4;
    wire OutReg_0_4_i_m3_ns_1_4_cascade_;
    wire OutReg_ess_RNO_1Z0Z_4;
    wire OutReg_0_5_i_m3_ns_1_4;
    wire ch0_A_c;
    wire \QuadInstance3.Quad_RNO_0_3_6 ;
    wire \QuadInstance6.Quad_RNO_0_6_4 ;
    wire dataRead6_4;
    wire \QuadInstance7.Quad_RNO_0_7_4 ;
    wire dataRead7_4;
    wire bfn_13_6_0_;
    wire \QuadInstance1.Quad_RNO_0_0_1 ;
    wire \QuadInstance1.un1_Quad_cry_0 ;
    wire \QuadInstance1.Quad_RNO_0_1_2 ;
    wire \QuadInstance1.un1_Quad_cry_1 ;
    wire \QuadInstance1.Quad_RNO_0_1_3 ;
    wire \QuadInstance1.un1_Quad_cry_2 ;
    wire \QuadInstance1.Quad_RNO_0_1_4 ;
    wire \QuadInstance1.un1_Quad_cry_3 ;
    wire \QuadInstance1.Quad_RNO_0_1_5 ;
    wire \QuadInstance1.un1_Quad_cry_4 ;
    wire \QuadInstance1.Quad_RNO_0_1_6 ;
    wire \QuadInstance1.un1_Quad_cry_5 ;
    wire \QuadInstance1.Quad_RNO_0_1_7 ;
    wire \QuadInstance1.un1_Quad_cry_6 ;
    wire \QuadInstance1.un1_Quad_cry_7 ;
    wire \QuadInstance1.Quad_RNO_0_1_8 ;
    wire bfn_13_7_0_;
    wire \QuadInstance1.un1_Quad_cry_8 ;
    wire \QuadInstance1.Quad_RNO_0_1_10 ;
    wire \QuadInstance1.un1_Quad_cry_9 ;
    wire \QuadInstance1.Quad_RNO_0_1_11 ;
    wire \QuadInstance1.un1_Quad_cry_10 ;
    wire \QuadInstance1.un1_Quad_cry_11 ;
    wire \QuadInstance1.un1_Quad_cry_12 ;
    wire \QuadInstance1.Quad_RNO_0_1_14 ;
    wire \QuadInstance1.un1_Quad_cry_13 ;
    wire \QuadInstance1.un1_Quad_cry_14 ;
    wire \QuadInstance6.Quad_RNO_0_6_9 ;
    wire \QuadInstance2.Quad_RNO_0_1_1 ;
    wire quadWriteZ0Z_2;
    wire \QuadInstance3.Quad_RNO_0_2_1 ;
    wire quadWriteZ0Z_3;
    wire \QuadInstance3.Quad_RNO_0_3_4 ;
    wire dataRead3_4;
    wire \QuadInstance1.Quad_RNO_0_1_9 ;
    wire \QuadInstance7.count_enable ;
    wire \QuadInstance6.delayedCh_BZ0Z_2 ;
    wire \QuadInstance6.Quad_RNIGENB1Z0Z_10 ;
    wire \QuadInstance6.delayedCh_AZ0Z_1 ;
    wire \QuadInstance6.delayedCh_AZ0Z_2 ;
    wire dataRead6_13;
    wire quadWriteZ0Z_6;
    wire \QuadInstance6.un1_count_enable_i_a2_0_1 ;
    wire \QuadInstance6.count_enable ;
    wire \QuadInstance6.Quad_RNIJHNB1Z0Z_13 ;
    wire \QuadInstance6.delayedCh_BZ0Z_1 ;
    wire dataRead2_11;
    wire dataRead3_11;
    wire OutReg_0_4_i_m3_i_m3_ns_1_11;
    wire dataRead5_12;
    wire dataRead2_12;
    wire dataRead3_12;
    wire dataRead6_12;
    wire dataRead7_12;
    wire OutReg_0_4_i_m3_ns_1_12_cascade_;
    wire OutReg_esr_RNO_1Z0Z_12_cascade_;
    wire OutReg_esr_RNO_2Z0Z_12;
    wire OutRegZ0Z_11;
    wire OutReg_esr_RNO_0Z0Z_12_cascade_;
    wire OutRegZ0Z_12;
    wire data_receivedZ0Z_12;
    wire data_receivedZ0Z_13;
    wire data_receivedZ0Z_14;
    wire data_receivedZ0Z_10;
    wire data_receivedZ0Z_11;
    wire data_received_esr_RNIMIH31Z0Z_19_cascade_;
    wire data_receivedZ0Z_19;
    wire data_receivedZ0Z_23;
    wire data_received_esr_RNIMIH31_0Z0Z_19_cascade_;
    wire \PWMInstance6.PWMPulseWidthCountZ0Z_5 ;
    wire \PWMInstance6.PWMPulseWidthCountZ0Z_8 ;
    wire \PWMInstance6.periodCounterZ0Z_15 ;
    wire \PWMInstance6.periodCounterZ0Z_14 ;
    wire \PWMInstance6.un1_PWMPulseWidthCount_0_I_21_c_RNO_5 ;
    wire \PWMInstance6.PWMPulseWidthCountZ0Z_14 ;
    wire \PWMInstance6.PWMPulseWidthCountZ0Z_15 ;
    wire \PWMInstance6.periodCounterZ0Z_10 ;
    wire \PWMInstance6.PWMPulseWidthCountZ0Z_11 ;
    wire \PWMInstance6.periodCounterZ0Z_11 ;
    wire \PWMInstance6.un1_PWMPulseWidthCount_0_I_33_c_RNO_5 ;
    wire \PWMInstance6.PWMPulseWidthCountZ0Z_10 ;
    wire \PWMInstance6.PWMPulseWidthCountZ0Z_13 ;
    wire \PWMInstance6.periodCounterZ0Z_12 ;
    wire \PWMInstance6.periodCounterZ0Z_13 ;
    wire \PWMInstance6.PWMPulseWidthCountZ0Z_12 ;
    wire \PWMInstance6.un1_PWMPulseWidthCount_0_I_39_c_RNO_5 ;
    wire \PWMInstance4.un1_periodCounter12_1_0_a2_0_0_cascade_ ;
    wire \PWMInstance4.PWMPulseWidthCountZ0Z_4 ;
    wire \PWMInstance4.PWMPulseWidthCountZ0Z_5 ;
    wire \PWMInstance4.PWMPulseWidthCountZ0Z_10 ;
    wire \PWMInstance4.PWMPulseWidthCountZ0Z_11 ;
    wire ch2_B_c;
    wire \QuadInstance2.delayedCh_BZ0Z_0 ;
    wire ch4_B_c;
    wire ch4_A_c;
    wire dataRead1_4;
    wire \QuadInstance1.Quad_RNIRK0OZ0Z_4 ;
    wire \QuadInstance1.delayedCh_BZ0Z_1 ;
    wire \QuadInstance1.count_enable_cascade_ ;
    wire \QuadInstance1.Quad_RNIOH0OZ0Z_1 ;
    wire \QuadInstance1.Quad_RNITM0OZ0Z_6 ;
    wire \QuadInstance1.Quad_RNISL0OZ0Z_5 ;
    wire \QuadInstance1.delayedCh_AZ0Z_2 ;
    wire \QuadInstance1.delayedCh_BZ0Z_2 ;
    wire \QuadInstance1.delayedCh_AZ0Z_1 ;
    wire \QuadInstance1.Quad_RNI0Q0OZ0Z_9 ;
    wire \QuadInstance1.Quad_RNI8P5DZ0Z_10 ;
    wire data_received_esr_RNIMIH31Z0Z_19;
    wire dataRead1_11;
    wire \QuadInstance1.Quad_RNI9Q5DZ0Z_11 ;
    wire dataRead3_5;
    wire dataRead2_5;
    wire \QuadInstance1.Quad_RNIUN0OZ0Z_7 ;
    wire \QuadInstance1.Quad_RNIPI0OZ0Z_2 ;
    wire \QuadInstance1.Quad_RNIQJ0OZ0Z_3 ;
    wire \QuadInstance1.Quad_RNIAR5DZ0Z_12 ;
    wire \QuadInstance1.Quad_RNIBS5DZ0Z_13 ;
    wire \QuadInstance1.Quad_RNICT5DZ0Z_14 ;
    wire \QuadInstance1.Quad_RNIVO0OZ0Z_8 ;
    wire \QuadInstance1.un1_count_enable_i_a2_0_1 ;
    wire \QuadInstance1.un1_Quad_axb_15 ;
    wire \QuadInstance1.count_enable ;
    wire \QuadInstance1.Quad_RNO_0_1_12 ;
    wire dataRead1_12;
    wire quadWriteZ0Z_1;
    wire \QuadInstance1.Quad_RNO_0_1_13 ;
    wire dataRead1_13;
    wire dataRead1_1;
    wire dataRead5_1;
    wire OutReg_ess_RNO_2Z0Z_1_cascade_;
    wire dataRead2_1;
    wire dataRead3_1;
    wire dataRead6_1;
    wire OutReg_0_4_i_m3_ns_1_1_cascade_;
    wire OutReg_ess_RNO_1Z0Z_1;
    wire OutReg_0_5_i_m3_ns_1_1;
    wire dataRead2_3;
    wire dataRead3_3;
    wire dataRead3_15;
    wire dataRead2_15;
    wire dataRead7_15;
    wire dataRead6_15;
    wire OutReg_0_4_i_m3_ns_1_15_cascade_;
    wire dataRead5_15;
    wire dataRead1_15;
    wire data_receivedZ0Z_5;
    wire data_receivedZ0Z_6;
    wire data_receivedZ0Z_7;
    wire data_receivedZ0Z_8;
    wire data_receivedZ0Z_9;
    wire N_870_i;
    wire pwmWriteZ0Z_3;
    wire pwmWrite_fastZ0Z_3;
    wire \PWMInstance3.clkCountZ0Z_1 ;
    wire \PWMInstance3.clkCountZ0Z_0 ;
    wire \PWMInstance3.un1_periodCounter12_1_0_a2_0_6_cascade_ ;
    wire \PWMInstance3.un1_periodCounter12_1_0_a2_0_14_cascade_ ;
    wire \PWMInstance6.PWMPulseWidthCountZ0Z_9 ;
    wire \PWMInstance6.pwmWrite_0_6 ;
    wire \PWMInstance4.PWMPulseWidthCountZ0Z_3 ;
    wire \PWMInstance4.PWMPulseWidthCountZ0Z_2 ;
    wire \PWMInstance4.PWMPulseWidthCountZ0Z_14 ;
    wire \PWMInstance4.PWMPulseWidthCountZ0Z_15 ;
    wire \PWMInstance4.PWMPulseWidthCountZ0Z_12 ;
    wire \PWMInstance4.PWMPulseWidthCountZ0Z_13 ;
    wire bfn_14_16_0_;
    wire \PWMInstance4.un1_periodCounter_2_cry_0 ;
    wire \PWMInstance4.periodCounterZ0Z_2 ;
    wire \PWMInstance4.un1_periodCounter_2_cry_1 ;
    wire \PWMInstance4.periodCounterZ0Z_3 ;
    wire \PWMInstance4.un1_periodCounter_2_cry_2 ;
    wire \PWMInstance4.periodCounterZ0Z_4 ;
    wire \PWMInstance4.un1_periodCounter_2_cry_3 ;
    wire \PWMInstance4.periodCounterZ0Z_5 ;
    wire \PWMInstance4.un1_periodCounter_2_cry_4 ;
    wire \PWMInstance4.un1_periodCounter_2_cry_5 ;
    wire \PWMInstance4.un1_periodCounter_2_cry_6 ;
    wire \PWMInstance4.un1_periodCounter_2_cry_7 ;
    wire bfn_14_17_0_;
    wire \PWMInstance4.un1_periodCounter_2_cry_8 ;
    wire \PWMInstance4.periodCounterZ0Z_10 ;
    wire \PWMInstance4.un1_periodCounter_2_cry_9 ;
    wire \PWMInstance4.periodCounterZ0Z_11 ;
    wire \PWMInstance4.un1_periodCounter_2_cry_10 ;
    wire \PWMInstance4.periodCounterZ0Z_12 ;
    wire \PWMInstance4.un1_periodCounter_2_cry_11 ;
    wire \PWMInstance4.un1_periodCounter_2_cry_12 ;
    wire \PWMInstance4.periodCounterZ0Z_14 ;
    wire \PWMInstance4.un1_periodCounter_2_cry_13 ;
    wire \PWMInstance4.un1_periodCounter_2_cry_14 ;
    wire \PWMInstance4.un1_periodCounter_2_cry_15 ;
    wire bfn_14_18_0_;
    wire bfn_15_1_0_;
    wire \PWMInstance4.un1_PWMPulseWidthCount_0_I_9_c_RNO_3 ;
    wire \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_0 ;
    wire \PWMInstance4.un1_PWMPulseWidthCount_0_I_15_c_RNO_3 ;
    wire \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_1 ;
    wire \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_2 ;
    wire \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_3 ;
    wire \PWMInstance4.un1_PWMPulseWidthCount_0_I_33_c_RNO_3 ;
    wire \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_4 ;
    wire \PWMInstance4.un1_PWMPulseWidthCount_0_I_39_c_RNO_3 ;
    wire \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_5 ;
    wire \PWMInstance4.un1_PWMPulseWidthCount_0_I_21_c_RNO_3 ;
    wire \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_6 ;
    wire \PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_7 ;
    wire bfn_15_2_0_;
    wire PWM4_c;
    wire bfn_15_3_0_;
    wire \QuadInstance4.Quad_RNO_0_3_1 ;
    wire \QuadInstance4.un1_Quad_cry_0 ;
    wire \QuadInstance4.un1_Quad_cry_1 ;
    wire \QuadInstance4.un1_Quad_cry_2 ;
    wire \QuadInstance4.Quad_RNO_0_4_4 ;
    wire \QuadInstance4.un1_Quad_cry_3 ;
    wire \QuadInstance4.un1_Quad_cry_4 ;
    wire \QuadInstance4.un1_Quad_cry_5 ;
    wire \QuadInstance4.un1_Quad_cry_6 ;
    wire \QuadInstance4.un1_Quad_cry_7 ;
    wire bfn_15_4_0_;
    wire \QuadInstance4.Quad_RNO_0_4_9 ;
    wire \QuadInstance4.un1_Quad_cry_8 ;
    wire \QuadInstance4.un1_Quad_cry_9 ;
    wire \QuadInstance4.un1_Quad_cry_10 ;
    wire \QuadInstance4.un1_Quad_cry_11 ;
    wire \QuadInstance4.un1_Quad_cry_12 ;
    wire \QuadInstance4.un1_Quad_cry_13 ;
    wire \QuadInstance4.un1_Quad_axb_15 ;
    wire \QuadInstance4.un1_Quad_cry_14 ;
    wire \QuadInstance4.Quad_RNO_0_4_6 ;
    wire \QuadInstance4.Quad_RNIL00S1Z0Z_6 ;
    wire \QuadInstance4.Quad_RNI06TL1Z0Z_10 ;
    wire \QuadInstance4.Quad_RNI17TL1Z0Z_11 ;
    wire \QuadInstance4.Quad_RNO_0_4_11 ;
    wire dataRead4_11;
    wire dataRead4_6;
    wire dataRead1_6;
    wire dataRead5_6;
    wire OutReg_0_5_i_m3_ns_1_6_cascade_;
    wire \QuadInstance4.Quad_RNIO30S1Z0Z_9 ;
    wire \QuadInstance4.Quad_RNIM10S1Z0Z_7 ;
    wire dataRead4_15;
    wire OutReg_0_5_i_m3_ns_1_15;
    wire dataRead1_9;
    wire dataRead5_9;
    wire OutReg_ess_RNO_2Z0Z_9_cascade_;
    wire dataRead3_9;
    wire dataRead2_9;
    wire dataRead6_9;
    wire dataRead7_9;
    wire OutReg_0_4_i_m3_ns_1_9_cascade_;
    wire OutReg_ess_RNO_1Z0Z_9;
    wire dataRead4_9;
    wire OutReg_0_5_i_m3_ns_1_9;
    wire N_45_0_g;
    wire N_1187_g;
    wire \QuadInstance4.Quad_RNO_0_4_13 ;
    wire \QuadInstance7.Quad_RNO_0_7_13 ;
    wire dataRead7_13;
    wire \QuadInstance4.Quad_RNO_0_4_3 ;
    wire \QuadInstance7.Quad_RNO_0_7_3 ;
    wire quadWriteZ0Z_7;
    wire \QuadInstance7.Quad_RNO_0_6_1 ;
    wire dataRead7_1;
    wire quadWriteZ0Z_5;
    wire \QuadInstance5.Quad_RNO_0_5_3 ;
    wire GB_BUFFER_RST_c_i_g_THRU_CO;
    wire dataRead5_7;
    wire dataRead1_7;
    wire OutReg_ess_RNO_2Z0Z_7_cascade_;
    wire OutReg_ess_RNO_0Z0Z_7_cascade_;
    wire dataRead2_7;
    wire dataRead3_7;
    wire dataRead6_7;
    wire dataRead7_7;
    wire OutReg_0_4_i_m3_ns_1_7_cascade_;
    wire OutReg_ess_RNO_1Z0Z_7;
    wire OutReg_ess_RNO_0Z0Z_9;
    wire OutRegZ0Z_13;
    wire OutRegZ0Z_14;
    wire \PWMInstance3.PWMPulseWidthCountZ0Z_5 ;
    wire \PWMInstance3.un1_periodCounter12_1_0_a2_0_0_cascade_ ;
    wire \PWMInstance3.un1_periodCounter12_1_0_a2_0_12 ;
    wire \PWMInstance3.PWMPulseWidthCountZ0Z_4 ;
    wire \PWMInstance3.PWMPulseWidthCountZ0Z_11 ;
    wire \PWMInstance3.PWMPulseWidthCountZ0Z_10 ;
    wire \PWMInstance3.periodCounter12 ;
    wire bfn_15_13_0_;
    wire \PWMInstance3.un1_periodCounter_2_cry_0 ;
    wire \PWMInstance3.un1_periodCounter_2_cry_1 ;
    wire \PWMInstance3.un1_periodCounter_2_cry_2 ;
    wire \PWMInstance3.periodCounterZ0Z_4 ;
    wire \PWMInstance3.un1_periodCounter_2_cry_3 ;
    wire \PWMInstance3.un1_periodCounter_2_cry_4 ;
    wire \PWMInstance3.un1_periodCounter_2_cry_5 ;
    wire \PWMInstance3.un1_periodCounter_2_cry_6 ;
    wire \PWMInstance3.un1_periodCounter_2_cry_7 ;
    wire bfn_15_14_0_;
    wire \PWMInstance3.un1_periodCounter_2_cry_8 ;
    wire \PWMInstance3.periodCounterZ0Z_10 ;
    wire \PWMInstance3.un1_periodCounter_2_cry_9 ;
    wire \PWMInstance3.un1_periodCounter_2_cry_10 ;
    wire \PWMInstance3.un1_periodCounter_2_cry_11 ;
    wire \PWMInstance3.un1_periodCounter_2_cry_12 ;
    wire \PWMInstance3.un1_periodCounter_2_cry_13 ;
    wire \PWMInstance3.un1_periodCounter_2_cry_14 ;
    wire \PWMInstance3.un1_periodCounter_2_cry_15 ;
    wire bfn_15_15_0_;
    wire \PWMInstance3.periodCounterZ0Z_16 ;
    wire \PWMInstance4.periodCounterZ0Z_13 ;
    wire \PWMInstance4.periodCounterZ0Z_0 ;
    wire \PWMInstance4.PWMPulseWidthCountZ0Z_0 ;
    wire \PWMInstance4.un1_PWMPulseWidthCount_0_I_1_c_RNO_3 ;
    wire \PWMInstance4.PWMPulseWidthCountZ0Z_1 ;
    wire \PWMInstance4.periodCounterZ0Z_6 ;
    wire \PWMInstance4.un1_PWMPulseWidthCount_0_I_27_c_RNO_3 ;
    wire \PWMInstance4.PWMPulseWidthCountZ0Z_6 ;
    wire \PWMInstance4.PWMPulseWidthCountZ0Z_7 ;
    wire \PWMInstance4.PWMPulseWidthCountZ0Z_9 ;
    wire \PWMInstance4.periodCounterZ0Z_8 ;
    wire \PWMInstance4.periodCounterZ0Z_9 ;
    wire \PWMInstance4.PWMPulseWidthCountZ0Z_8 ;
    wire \PWMInstance4.un1_PWMPulseWidthCount_0_I_45_c_RNO_3 ;
    wire \PWMInstance4.un1_periodCounter12_1_0_a2_0 ;
    wire \PWMInstance4.periodCounterZ0Z_16 ;
    wire \PWMInstance4.periodCounterZ0Z_7 ;
    wire pwmWriteZ0Z_4;
    wire \PWMInstance4.pwmWrite_0_4 ;
    wire pwmWrite_fastZ0Z_4;
    wire \PWMInstance4.clkCountZ0Z_1 ;
    wire \PWMInstance4.clkCountZ0Z_0 ;
    wire \PWMInstance4.periodCounter12 ;
    wire \PWMInstance4.periodCounterZ0Z_15 ;
    wire \PWMInstance4.periodCounterZ0Z_1 ;
    wire \PWMInstance4.periodCounter12_cascade_ ;
    wire \PWMInstance4.un1_periodCounter12_1_0_a2_0_6 ;
    wire \PWMInstance4.un1_periodCounter12_1_0_a2_0_10 ;
    wire \PWMInstance4.un1_periodCounter12_1_0_a2_0_9 ;
    wire \PWMInstance4.un1_periodCounter12_1_0_a2_0_14_cascade_ ;
    wire \PWMInstance4.un1_periodCounter12_1_0_a2_0_12 ;
    wire \PWMInstance4.out_0_sqmuxa ;
    wire ch6_B_c;
    wire \QuadInstance6.delayedCh_BZ0Z_0 ;
    wire PWM4_obufLegalizeSB_DFFNet;
    wire ch1_B_c;
    wire \QuadInstance1.delayedCh_BZ0Z_0 ;
    wire \QuadInstance4.Quad_RNO_0_4_5 ;
    wire dataRead4_5;
    wire \QuadInstance4.Quad_RNIKVVR1Z0Z_5 ;
    wire \QuadInstance4.Quad_RNI28TL1Z0Z_12 ;
    wire \QuadInstance4.count_enable_cascade_ ;
    wire \QuadInstance4.Quad_RNIHSVR1Z0Z_2 ;
    wire dataRead4_1;
    wire \QuadInstance4.Quad_RNIGRVR1Z0Z_1 ;
    wire \QuadInstance4.Quad_RNO_0_4_2 ;
    wire dataRead4_2;
    wire \QuadInstance4.Quad_RNIITVR1Z0Z_3 ;
    wire \QuadInstance4.Quad_RNI39TL1Z0Z_13 ;
    wire \QuadInstance4.Quad_RNI4ATL1Z0Z_14 ;
    wire \QuadInstance4.delayedCh_BZ0Z_2 ;
    wire dataRead4_4;
    wire \QuadInstance4.un1_count_enable_i_a2_0_1_cascade_ ;
    wire \QuadInstance4.Quad_RNIJUVR1Z0Z_4 ;
    wire \QuadInstance4.delayedCh_AZ0Z_0 ;
    wire \QuadInstance4.delayedCh_AZ0Z_1 ;
    wire \QuadInstance4.delayedCh_AZ0Z_2 ;
    wire \QuadInstance4.count_enable ;
    wire \QuadInstance4.un1_count_enable_i_a2_0_1 ;
    wire \QuadInstance4.Quad_RNIN20S1Z0Z_8 ;
    wire \QuadInstance4.Quad_RNO_0_4_8 ;
    wire dataRead4_8;
    wire OutReg_0_5_i_m3_ns_1_7;
    wire \QuadInstance4.Quad_RNO_0_4_7 ;
    wire dataRead4_7;
    wire OutReg_0_5_i_m3_ns_1_12;
    wire \QuadInstance4.Quad_RNO_0_4_12 ;
    wire dataRead4_12;
    wire dataRead4_13;
    wire OutReg_0_5_i_m3_ns_1_13;
    wire data_received_2_repZ0Z1;
    wire dataRead4_3;
    wire data_received_0_repZ0Z1;
    wire dataRead5_3;
    wire dataRead1_3;
    wire OutReg_0_5_i_m3_ns_1_3_cascade_;
    wire dataRead7_3;
    wire dataRead6_3;
    wire OutReg_0_4_i_m3_ns_1_3;
    wire OutReg_ess_RNO_1Z0Z_3_cascade_;
    wire OutReg_ess_RNO_2Z0Z_3;
    wire OutReg_ess_RNO_0Z0Z_3_cascade_;
    wire OutRegZ0Z_3;
    wire OutReg_ess_RNO_0Z0Z_4;
    wire dataRead6_6;
    wire dataRead7_6;
    wire OutReg_esr_RNO_1Z0Z_6_cascade_;
    wire OutReg_esr_RNO_2Z0Z_6;
    wire OutReg_esr_RNO_0Z0Z_6_cascade_;
    wire OutRegZ0Z_6;
    wire dataRead2_6;
    wire dataRead3_6;
    wire OutReg_0_4_i_m3_ns_1_6;
    wire dataRead5_14;
    wire dataRead1_14;
    wire OutReg_0_5_i_m3_ns_1_14_cascade_;
    wire OutReg_esr_RNO_2Z0Z_14_cascade_;
    wire OutReg_esr_RNO_1Z0Z_14;
    wire OutReg_esr_RNO_0Z0Z_14;
    wire dataWriteZ0Z_8;
    wire dataWriteZ0Z_12;
    wire dataWriteZ0Z_13;
    wire dataWriteZ0Z_9;
    wire \PWMInstance3.periodCounterZ0Z_5 ;
    wire \PWMInstance3.periodCounterZ0Z_11 ;
    wire \PWMInstance3.un1_periodCounter12_1_0_a2_0_10 ;
    wire \PWMInstance3.PWMPulseWidthCountZ0Z_3 ;
    wire \PWMInstance3.periodCounterZ0Z_3 ;
    wire \PWMInstance3.periodCounterZ0Z_2 ;
    wire \PWMInstance3.PWMPulseWidthCountZ0Z_2 ;
    wire \PWMInstance3.periodCounterZ0Z_15 ;
    wire \PWMInstance3.periodCounterZ0Z_14 ;
    wire \PWMInstance3.PWMPulseWidthCountZ0Z_14 ;
    wire \PWMInstance3.PWMPulseWidthCountZ0Z_15 ;
    wire \PWMInstance3.PWMPulseWidthCountZ0Z_13 ;
    wire \PWMInstance3.PWMPulseWidthCountZ0Z_12 ;
    wire \PWMInstance3.periodCounterZ0Z_12 ;
    wire \PWMInstance3.periodCounterZ0Z_13 ;
    wire \PWMInstance3.un1_periodCounter12_1_0_a2_0_9 ;
    wire \PWMInstance3.periodCounterZ0Z_0 ;
    wire \PWMInstance3.periodCounterZ0Z_1 ;
    wire \PWMInstance3.PWMPulseWidthCountZ0Z_0 ;
    wire \PWMInstance3.PWMPulseWidthCountZ0Z_1 ;
    wire \PWMInstance3.periodCounterZ0Z_7 ;
    wire \PWMInstance3.periodCounterZ0Z_6 ;
    wire \PWMInstance3.PWMPulseWidthCountZ0Z_6 ;
    wire dataWriteZ0Z_7;
    wire \PWMInstance3.PWMPulseWidthCountZ0Z_7 ;
    wire \PWMInstance3.pwmWrite_0_3 ;
    wire \PWMInstance3.PWMPulseWidthCountZ0Z_8 ;
    wire \PWMInstance3.periodCounterZ0Z_8 ;
    wire \PWMInstance3.periodCounterZ0Z_9 ;
    wire \PWMInstance3.PWMPulseWidthCountZ0Z_9 ;
    wire \PWMInstance3.un1_PWMPulseWidthCount_0_I_1_c_RNO_2 ;
    wire bfn_16_15_0_;
    wire \PWMInstance3.un1_PWMPulseWidthCount_0_I_9_c_RNO_2 ;
    wire \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_0 ;
    wire \PWMInstance3.un1_PWMPulseWidthCount_0_I_15_c_RNO_2 ;
    wire \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_1 ;
    wire \PWMInstance3.un1_PWMPulseWidthCount_0_I_27_c_RNO_2 ;
    wire \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_2 ;
    wire \PWMInstance3.un1_PWMPulseWidthCount_0_I_45_c_RNO_2 ;
    wire \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_3 ;
    wire \PWMInstance3.un1_PWMPulseWidthCount_0_I_33_c_RNO_2 ;
    wire \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_4 ;
    wire \PWMInstance3.un1_PWMPulseWidthCount_0_I_39_c_RNO_2 ;
    wire \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_5 ;
    wire \PWMInstance3.un1_PWMPulseWidthCount_0_I_21_c_RNO_2 ;
    wire \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_6 ;
    wire \PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_7 ;
    wire \PWMInstance3.un1_periodCounter12_1_0_a2_0 ;
    wire \PWMInstance3.out_0_sqmuxa ;
    wire bfn_16_16_0_;
    wire PWM3_c;
    wire ch7_A_c;
    wire \QuadInstance7.delayedCh_AZ0Z_0 ;
    wire \QuadInstance4.Quad_RNO_0_4_10 ;
    wire quadWriteZ0Z_4;
    wire \QuadInstance4.Quad_RNO_0_4_14 ;
    wire dataRead4_14;
    wire \QuadInstance0.delayedCh_BZ0Z_0 ;
    wire \QuadInstance4.delayedCh_BZ0Z_0 ;
    wire \QuadInstance4.delayedCh_BZ0Z_1 ;
    wire bfn_17_6_0_;
    wire \QuadInstance0.Quad_RNO_0Z0Z_1 ;
    wire \QuadInstance0.un1_Quad_cry_0 ;
    wire \QuadInstance0.Quad_RNO_0_0_2 ;
    wire \QuadInstance0.un1_Quad_cry_1 ;
    wire \QuadInstance0.Quad_RNO_0_0_3 ;
    wire \QuadInstance0.un1_Quad_cry_2 ;
    wire \QuadInstance0.Quad_RNO_0_0_4 ;
    wire \QuadInstance0.un1_Quad_cry_3 ;
    wire \QuadInstance0.Quad_RNO_0_0_5 ;
    wire \QuadInstance0.un1_Quad_cry_4 ;
    wire \QuadInstance0.Quad_RNO_0_0_6 ;
    wire \QuadInstance0.un1_Quad_cry_5 ;
    wire dataRead0_7;
    wire \QuadInstance0.Quad_RNIMKBH1Z0Z_7 ;
    wire \QuadInstance0.Quad_RNO_0_0_7 ;
    wire \QuadInstance0.un1_Quad_cry_6 ;
    wire \QuadInstance0.un1_Quad_cry_7 ;
    wire dataRead0_8;
    wire \QuadInstance0.Quad_RNINLBH1Z0Z_8 ;
    wire \QuadInstance0.Quad_RNO_0_0_8 ;
    wire bfn_17_7_0_;
    wire dataRead0_9;
    wire \QuadInstance0.Quad_RNIOMBH1Z0Z_9 ;
    wire \QuadInstance0.Quad_RNO_0_0_9 ;
    wire \QuadInstance0.un1_Quad_cry_8 ;
    wire \QuadInstance0.un1_Quad_cry_9 ;
    wire dataRead0_11;
    wire \QuadInstance0.Quad_RNI1M8Q1Z0Z_11 ;
    wire \QuadInstance0.Quad_RNO_0_0_11 ;
    wire \QuadInstance0.un1_Quad_cry_10 ;
    wire dataRead0_12;
    wire \QuadInstance0.Quad_RNI2N8Q1Z0Z_12 ;
    wire \QuadInstance0.Quad_RNO_0_0_12 ;
    wire \QuadInstance0.un1_Quad_cry_11 ;
    wire dataRead0_13;
    wire \QuadInstance0.Quad_RNI3O8Q1Z0Z_13 ;
    wire \QuadInstance0.Quad_RNO_0_0_13 ;
    wire \QuadInstance0.un1_Quad_cry_12 ;
    wire \QuadInstance0.un1_Quad_cry_13 ;
    wire \QuadInstance0.un1_Quad_axb_15 ;
    wire \QuadInstance0.un1_Quad_cry_14 ;
    wire dataRead0_15;
    wire dataRead1_2;
    wire dataRead5_2;
    wire OutReg_0_5_i_m3_ns_1_2;
    wire OutReg_esr_RNO_2Z0Z_2_cascade_;
    wire OutReg_esr_RNO_0Z0Z_2_cascade_;
    wire OutRegZ0Z_2;
    wire dataRead2_2;
    wire dataRead3_2;
    wire dataRead7_2;
    wire dataRead6_2;
    wire OutReg_0_4_i_m3_ns_1_2_cascade_;
    wire OutReg_esr_RNO_1Z0Z_2;
    wire dataRead0_0;
    wire dataRead4_0;
    wire dataRead1_0;
    wire OutReg_0_5_i_m3_ns_1_0_cascade_;
    wire dataRead5_0;
    wire OutReg_ess_RNO_1Z0Z_0_cascade_;
    wire dataRead3_0;
    wire dataRead2_0;
    wire dataRead6_0;
    wire OutReg_0_4_i_m3_ns_1_0_cascade_;
    wire dataRead7_0;
    wire OutReg_ess_RNO_0Z0Z_0;
    wire OutRegZ0Z_0;
    wire OutReg_ess_RNO_0Z0Z_1;
    wire OutRegZ0Z_1;
    wire dataRead2_8;
    wire dataRead3_8;
    wire data_receivedZ0Z_3;
    wire data_received_esr_RNI7L871Z0Z_3_cascade_;
    wire OutReg_0_sqmuxa_0_a2_3_a2_2;
    wire dataWriteZ0Z_0;
    wire \PWMInstance2.PWMPulseWidthCountZ0Z_0 ;
    wire dataWriteZ0Z_1;
    wire \PWMInstance2.PWMPulseWidthCountZ0Z_1 ;
    wire \PWMInstance2.PWMPulseWidthCountZ0Z_7 ;
    wire dataWriteZ0Z_6;
    wire \PWMInstance2.PWMPulseWidthCountZ0Z_6 ;
    wire \PWMInstance2.PWMPulseWidthCountZ0Z_8 ;
    wire \PWMInstance2.PWMPulseWidthCountZ0Z_9 ;
    wire pwmWriteZ0Z_2;
    wire pwmWrite_fastZ0Z_2;
    wire \PWMInstance2.clkCountZ0Z_1 ;
    wire \PWMInstance2.clkCountZ0Z_0 ;
    wire \PWMInstance2.un1_periodCounter12_1_0_a2_0_6_cascade_ ;
    wire \PWMInstance2.un1_periodCounter12_1_0_a2_0_9 ;
    wire \PWMInstance2.un1_periodCounter12_1_0_a2_0_14_cascade_ ;
    wire \PWMInstance2.un1_periodCounter12_1_0_a2_0_10 ;
    wire dataWriteZ0Z_2;
    wire \PWMInstance2.PWMPulseWidthCountZ0Z_2 ;
    wire dataWriteZ0Z_3;
    wire \PWMInstance2.PWMPulseWidthCountZ0Z_3 ;
    wire \PWMInstance2.PWMPulseWidthCountZ0Z_14 ;
    wire dataWriteZ0Z_15;
    wire \PWMInstance2.PWMPulseWidthCountZ0Z_15 ;
    wire \PWMInstance2.PWMPulseWidthCountZ0Z_13 ;
    wire \PWMInstance2.PWMPulseWidthCountZ0Z_12 ;
    wire \PWMInstance2.un1_PWMPulseWidthCount_0_I_1_c_RNO_1 ;
    wire bfn_17_14_0_;
    wire \PWMInstance2.un1_PWMPulseWidthCount_0_I_9_c_RNO_1 ;
    wire \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_0 ;
    wire \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_1 ;
    wire \PWMInstance2.un1_PWMPulseWidthCount_0_I_27_c_RNO_1 ;
    wire \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_2 ;
    wire \PWMInstance2.un1_PWMPulseWidthCount_0_I_45_c_RNO_1 ;
    wire \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_3 ;
    wire \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_4 ;
    wire \PWMInstance2.un1_PWMPulseWidthCount_0_I_39_c_RNO_1 ;
    wire \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_5 ;
    wire CONSTANT_ONE_NET;
    wire \PWMInstance2.un1_PWMPulseWidthCount_0_I_21_c_RNO_1 ;
    wire \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_6 ;
    wire \PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_7 ;
    wire \PWMInstance2.un1_periodCounter12_1_0_a2_0 ;
    wire bfn_17_15_0_;
    wire PWM2_c;
    wire MOSI_c;
    wire ch1_A_c;
    wire \QuadInstance1.delayedCh_AZ0Z_0 ;
    wire \QuadInstance0.delayedCh_AZ0Z_0 ;
    wire data_received_0_repZ0Z2;
    wire dataRead4_10;
    wire data_received_2_repZ0Z2;
    wire \QuadInstance0.Quad_RNO_0_0_10 ;
    wire \QuadInstance0.delayedCh_BZ0Z_1 ;
    wire \QuadInstance0.delayedCh_AZ0Z_2 ;
    wire dataRead0_1;
    wire \QuadInstance0.count_enable_cascade_ ;
    wire \QuadInstance0.Quad_RNIGEBH1Z0Z_1 ;
    wire dataRead0_10;
    wire \QuadInstance0.Quad_RNI0L8Q1Z0Z_10 ;
    wire dataRead0_2;
    wire \QuadInstance0.Quad_RNIHFBH1Z0Z_2 ;
    wire \QuadInstance0.delayedCh_BZ0Z_2 ;
    wire \QuadInstance0.delayedCh_AZ0Z_1 ;
    wire RST_c;
    wire dataWriteZ0Z_14;
    wire \QuadInstance0.Quad_RNO_0_0_14 ;
    wire dataRead0_14;
    wire \QuadInstance0.Quad_RNI4P8Q1Z0Z_14 ;
    wire dataRead0_3;
    wire \QuadInstance0.Quad_RNIIGBH1Z0Z_3 ;
    wire dataRead0_4;
    wire \QuadInstance0.Quad_RNIJHBH1Z0Z_4 ;
    wire dataRead0_5;
    wire \QuadInstance0.Quad_RNIKIBH1Z0Z_5 ;
    wire \QuadInstance0.count_enable ;
    wire dataRead0_6;
    wire \QuadInstance0.un1_count_enable_i_a2_0_1 ;
    wire \QuadInstance0.Quad_RNILJBH1Z0Z_6 ;
    wire data_receivedZ0Z_21;
    wire data_receivedZ0Z_20;
    wire data_receivedZ0Z_22;
    wire data_received_esr_RNIMIH31_0Z0Z_19;
    wire quadWriteZ0Z_0;
    wire MOSIrZ0Z_0;
    wire MOSIrZ0Z_1;
    wire dataRead1_10;
    wire dataRead5_10;
    wire OutReg_0_5_i_m3_ns_1_10;
    wire data_receivedZ0Z_4;
    wire un1_OutReg51_4_0_i_o3_2_cascade_;
    wire OutReg_21_m_0_a2_1_0;
    wire OutReg_esr_RNO_2Z0Z_10;
    wire OutRegZ0Z_9;
    wire OutReg_esr_RNO_0Z0Z_10;
    wire OutRegZ0Z_10;
    wire data_received_fastZ0Z_2;
    wire dataRead3_10;
    wire data_received_fastZ0Z_0;
    wire dataRead2_10;
    wire dataRead7_10;
    wire dataRead6_10;
    wire OutReg_0_4_i_m3_ns_1_10_cascade_;
    wire OutReg_esr_RNO_1Z0Z_10;
    wire \PWMInstance2.periodCounter12 ;
    wire \PWMInstance2.periodCounterZ0Z_0 ;
    wire bfn_18_11_0_;
    wire \PWMInstance2.periodCounterZ0Z_1 ;
    wire \PWMInstance2.un1_periodCounter_2_cry_0 ;
    wire \PWMInstance2.un1_periodCounter_2_cry_1 ;
    wire \PWMInstance2.periodCounterZ0Z_3 ;
    wire \PWMInstance2.un1_periodCounter_2_cry_2 ;
    wire \PWMInstance2.un1_periodCounter_2_cry_3 ;
    wire \PWMInstance2.un1_periodCounter_2_cry_4 ;
    wire \PWMInstance2.periodCounterZ0Z_6 ;
    wire \PWMInstance2.un1_periodCounter_2_cry_5 ;
    wire \PWMInstance2.periodCounterZ0Z_7 ;
    wire \PWMInstance2.un1_periodCounter_2_cry_6 ;
    wire \PWMInstance2.un1_periodCounter_2_cry_7 ;
    wire \PWMInstance2.periodCounterZ0Z_8 ;
    wire bfn_18_12_0_;
    wire \PWMInstance2.periodCounterZ0Z_9 ;
    wire \PWMInstance2.un1_periodCounter_2_cry_8 ;
    wire \PWMInstance2.un1_periodCounter_2_cry_9 ;
    wire \PWMInstance2.un1_periodCounter_2_cry_10 ;
    wire \PWMInstance2.un1_periodCounter_2_cry_11 ;
    wire \PWMInstance2.periodCounterZ0Z_13 ;
    wire \PWMInstance2.un1_periodCounter_2_cry_12 ;
    wire \PWMInstance2.un1_periodCounter_2_cry_13 ;
    wire \PWMInstance2.periodCounterZ0Z_15 ;
    wire \PWMInstance2.un1_periodCounter_2_cry_14 ;
    wire \PWMInstance2.un1_periodCounter_2_cry_15 ;
    wire \PWMInstance2.out_0_sqmuxa ;
    wire bfn_18_13_0_;
    wire \PWMInstance2.periodCounterZ0Z_16 ;
    wire PWMInstance0_N_42_g;
    wire \PWMInstance2.periodCounterZ0Z_5 ;
    wire \PWMInstance2.un1_PWMPulseWidthCount_0_I_15_c_RNO_1 ;
    wire \PWMInstance2.periodCounterZ0Z_14 ;
    wire \PWMInstance2.periodCounterZ0Z_2 ;
    wire \PWMInstance2.periodCounterZ0Z_4 ;
    wire \PWMInstance2.periodCounterZ0Z_12 ;
    wire \PWMInstance2.un1_periodCounter12_1_0_a2_0_0_cascade_ ;
    wire \PWMInstance2.un1_periodCounter12_1_0_a2_0_12 ;
    wire dataWriteZ0Z_4;
    wire \PWMInstance2.PWMPulseWidthCountZ0Z_4 ;
    wire dataWriteZ0Z_5;
    wire \PWMInstance2.PWMPulseWidthCountZ0Z_5 ;
    wire \PWMInstance2.periodCounterZ0Z_10 ;
    wire \PWMInstance2.periodCounterZ0Z_11 ;
    wire \PWMInstance2.un1_PWMPulseWidthCount_0_I_33_c_RNO_1 ;
    wire dataWriteZ0Z_10;
    wire \PWMInstance2.PWMPulseWidthCountZ0Z_10 ;
    wire dataWriteZ0Z_11;
    wire \PWMInstance2.PWMPulseWidthCountZ0Z_11 ;
    wire \PWMInstance2.pwmWrite_0_2 ;
    wire RST_c_i_g;
    wire PWM2_obufLegalizeSB_DFFNet;
    wire PWM3_obufLegalizeSB_DFFNet;
    wire MISO_obufLegalizeSB_DFFNet;
    wire internalOscilatorOutputNet;
    wire dataRead5_5;
    wire dataRead1_5;
    wire OutReg_0_5_i_m3_ns_1_5;
    wire dataRead6_5;
    wire dataRead7_5;
    wire OutReg_0_4_i_m3_ns_1_5;
    wire OutReg_ess_RNO_1Z0Z_5_cascade_;
    wire OutReg_ess_RNO_2Z0Z_5;
    wire OutReg_ess_RNO_0Z0Z_5;
    wire OutRegZ0Z_4;
    wire OutRegZ0Z_5;
    wire OutRegZ0Z_15;
    wire dataOut_RNOZ0Z_0_cascade_;
    wire MISO_c;
    wire SSEL_c;
    wire un1_bit_count_1_c1_cascade_;
    wire OutReg_ess_RNO_1Z0Z_15;
    wire OutReg_ess_RNO_2Z0Z_15;
    wire OutReg_ess_RNO_0Z0Z_15;
    wire bit_countZ0Z_0;
    wire dataRead6_8;
    wire data_receivedZ0Z_2;
    wire dataRead7_8;
    wire OutReg_0_4_i_m3_ns_1_8;
    wire data_receivedZ0Z_1;
    wire OutReg_esr_RNO_1Z0Z_8_cascade_;
    wire OutRegZ0Z_7;
    wire OutReg_esr_RNO_0Z0Z_8_cascade_;
    wire un1_OutReg51_4_0_i_o3_2;
    wire OutRegZ0Z_8;
    wire N_863_0;
    wire OutReg_0_sqmuxa;
    wire dataRead1_8;
    wire dataRead5_8;
    wire data_receivedZ0Z_0;
    wire OutReg_0_5_i_m3_ns_1_8;
    wire OutReg_esr_RNO_2Z0Z_8;
    wire SSELrZ0Z_0;
    wire SSELrZ0Z_2;
    wire SCK_c;
    wire bit_countZ0Z_2;
    wire SCKr_RNIBA7CZ0Z_2;
    wire SCKr_RNIBA7CZ0Z_2_cascade_;
    wire N_45_0;
    wire SCKrZ0Z_0;
    wire un1_bit_count_1_c1;
    wire bit_countZ0Z_1;
    wire bit_count_RNIU615_0Z0Z_4;
    wire bit_count_RNIU615_0Z0Z_4_cascade_;
    wire SSELr_RNIGO0FZ0Z_1;
    wire SSELrZ0Z_1;
    wire un1_bit_count_1_c3;
    wire bit_countZ0Z_3;
    wire bit_countZ0Z_4;
    wire un1_OutReg51_4_0_i_o3_3;
    wire SCKrZ0Z_1;
    wire SCKrZ0Z_2;
    wire myclk;
    wire _gnd_net_;

    IO_PAD CLK_ibuf_iopad (
            .OE(N__39370),
            .DIN(N__39369),
            .DOUT(N__39368),
            .PACKAGEPIN(CLK));
    defparam CLK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK_ibuf_preio (
            .PADOEN(N__39370),
            .PADOUT(N__39369),
            .PADIN(N__39368),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PWM5_obuf_iopad (
            .OE(N__39361),
            .DIN(N__39360),
            .DOUT(N__39359),
            .PACKAGEPIN(PWM5));
    defparam PWM5_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PWM5_obuf_preio.PIN_TYPE=6'b101001;
    PRE_IO PWM5_obuf_preio (
            .PADOEN(N__39361),
            .PADOUT(N__39360),
            .PADIN(N__39359),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__21357),
            .DIN0(),
            .DOUT0(N__16401),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ch6_A_ibuf_iopad.PULLUP=1'b1;
    IO_PAD ch6_A_ibuf_iopad (
            .OE(N__39352),
            .DIN(N__39351),
            .DOUT(N__39350),
            .PACKAGEPIN(ch6_A));
    defparam ch6_A_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ch6_A_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ch6_A_ibuf_preio (
            .PADOEN(N__39352),
            .PADOUT(N__39351),
            .PADIN(N__39350),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ch6_A_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ch6_B_ibuf_iopad.PULLUP=1'b1;
    IO_PAD ch6_B_ibuf_iopad (
            .OE(N__39343),
            .DIN(N__39342),
            .DOUT(N__39341),
            .PACKAGEPIN(ch6_B));
    defparam ch6_B_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ch6_B_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ch6_B_ibuf_preio (
            .PADOEN(N__39343),
            .PADOUT(N__39342),
            .PADIN(N__39341),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ch6_B_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ch5_B_ibuf_iopad.PULLUP=1'b1;
    IO_PAD ch5_B_ibuf_iopad (
            .OE(N__39334),
            .DIN(N__39333),
            .DOUT(N__39332),
            .PACKAGEPIN(ch5_B));
    defparam ch5_B_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ch5_B_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ch5_B_ibuf_preio (
            .PADOEN(N__39334),
            .PADOUT(N__39333),
            .PADIN(N__39332),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ch5_B_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ch0_B_ibuf_iopad.PULLUP=1'b1;
    IO_PAD ch0_B_ibuf_iopad (
            .OE(N__39325),
            .DIN(N__39324),
            .DOUT(N__39323),
            .PACKAGEPIN(ch0_B));
    defparam ch0_B_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ch0_B_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ch0_B_ibuf_preio (
            .PADOEN(N__39325),
            .PADOUT(N__39324),
            .PADIN(N__39323),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ch0_B_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PWM6_obuf_iopad (
            .OE(N__39316),
            .DIN(N__39315),
            .DOUT(N__39314),
            .PACKAGEPIN(PWM6));
    defparam PWM6_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PWM6_obuf_preio.PIN_TYPE=6'b101001;
    PRE_IO PWM6_obuf_preio (
            .PADOEN(N__39316),
            .PADOUT(N__39315),
            .PADIN(N__39314),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__17397),
            .DIN0(),
            .DOUT0(N__21378),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PWM4_obuf_iopad (
            .OE(N__39307),
            .DIN(N__39306),
            .DOUT(N__39305),
            .PACKAGEPIN(PWM4));
    defparam PWM4_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PWM4_obuf_preio.PIN_TYPE=6'b101001;
    PRE_IO PWM4_obuf_preio (
            .PADOEN(N__39307),
            .PADOUT(N__39306),
            .PADIN(N__39305),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__27090),
            .DIN0(),
            .DOUT0(N__24981),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam RST_ibuf_iopad.PULLUP=1'b1;
    IO_PAD RST_ibuf_iopad (
            .OE(N__39298),
            .DIN(N__39297),
            .DOUT(N__39296),
            .PACKAGEPIN(RST));
    defparam RST_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RST_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RST_ibuf_preio (
            .PADOEN(N__39298),
            .PADOUT(N__39297),
            .PADIN(N__39296),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RST_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MISO_obuf_iopad (
            .OE(N__39289),
            .DIN(N__39288),
            .DOUT(N__39287),
            .PACKAGEPIN(MISO));
    defparam MISO_obuf_preio.NEG_TRIGGER=1'b0;
    defparam MISO_obuf_preio.PIN_TYPE=6'b101001;
    PRE_IO MISO_obuf_preio (
            .PADOEN(N__39289),
            .PADOUT(N__39288),
            .PADIN(N__39287),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__36942),
            .DIN0(),
            .DOUT0(N__36639),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ch5_A_ibuf_iopad.PULLUP=1'b1;
    IO_PAD ch5_A_ibuf_iopad (
            .OE(N__39280),
            .DIN(N__39279),
            .DOUT(N__39278),
            .PACKAGEPIN(ch5_A));
    defparam ch5_A_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ch5_A_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ch5_A_ibuf_preio (
            .PADOEN(N__39280),
            .PADOUT(N__39279),
            .PADIN(N__39278),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ch5_A_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ch2_B_ibuf_iopad.PULLUP=1'b1;
    IO_PAD ch2_B_ibuf_iopad (
            .OE(N__39271),
            .DIN(N__39270),
            .DOUT(N__39269),
            .PACKAGEPIN(ch2_B));
    defparam ch2_B_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ch2_B_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ch2_B_ibuf_preio (
            .PADOEN(N__39271),
            .PADOUT(N__39270),
            .PADIN(N__39269),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ch2_B_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ch4_B_ibuf_iopad.PULLUP=1'b1;
    IO_PAD ch4_B_ibuf_iopad (
            .OE(N__39262),
            .DIN(N__39261),
            .DOUT(N__39260),
            .PACKAGEPIN(ch4_B));
    defparam ch4_B_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ch4_B_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ch4_B_ibuf_preio (
            .PADOEN(N__39262),
            .PADOUT(N__39261),
            .PADIN(N__39260),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ch4_B_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PWM3_obuf_iopad (
            .OE(N__39253),
            .DIN(N__39252),
            .DOUT(N__39251),
            .PACKAGEPIN(PWM3));
    defparam PWM3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PWM3_obuf_preio.PIN_TYPE=6'b101001;
    PRE_IO PWM3_obuf_preio (
            .PADOEN(N__39253),
            .PADOUT(N__39252),
            .PADIN(N__39251),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__36948),
            .DIN0(),
            .DOUT0(N__29727),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PWM1_obuf_iopad (
            .OE(N__39244),
            .DIN(N__39243),
            .DOUT(N__39242),
            .PACKAGEPIN(PWM1));
    defparam PWM1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PWM1_obuf_preio.PIN_TYPE=6'b101001;
    PRE_IO PWM1_obuf_preio (
            .PADOEN(N__39244),
            .PADOUT(N__39243),
            .PADIN(N__39242),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__17403),
            .DIN0(),
            .DOUT0(N__15735),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ch4_A_ibuf_iopad.PULLUP=1'b1;
    IO_PAD ch4_A_ibuf_iopad (
            .OE(N__39235),
            .DIN(N__39234),
            .DOUT(N__39233),
            .PACKAGEPIN(ch4_A));
    defparam ch4_A_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ch4_A_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ch4_A_ibuf_preio (
            .PADOEN(N__39235),
            .PADOUT(N__39234),
            .PADIN(N__39233),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ch4_A_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ch7_A_ibuf_iopad.PULLUP=1'b1;
    IO_PAD ch7_A_ibuf_iopad (
            .OE(N__39226),
            .DIN(N__39225),
            .DOUT(N__39224),
            .PACKAGEPIN(ch7_A));
    defparam ch7_A_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ch7_A_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ch7_A_ibuf_preio (
            .PADOEN(N__39226),
            .PADOUT(N__39225),
            .PADIN(N__39224),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ch7_A_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ch3_B_ibuf_iopad.PULLUP=1'b1;
    IO_PAD ch3_B_ibuf_iopad (
            .OE(N__39217),
            .DIN(N__39216),
            .DOUT(N__39215),
            .PACKAGEPIN(ch3_B));
    defparam ch3_B_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ch3_B_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ch3_B_ibuf_preio (
            .PADOEN(N__39217),
            .PADOUT(N__39216),
            .PADIN(N__39215),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ch3_B_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PWM7_obuf_iopad (
            .OE(N__39208),
            .DIN(N__39207),
            .DOUT(N__39206),
            .PACKAGEPIN(PWM7));
    defparam PWM7_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PWM7_obuf_preio.PIN_TYPE=6'b101001;
    PRE_IO PWM7_obuf_preio (
            .PADOEN(N__39208),
            .PADOUT(N__39207),
            .PADIN(N__39206),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__17391),
            .DIN0(),
            .DOUT0(N__14895),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SCK_ibuf_iopad (
            .OE(N__39199),
            .DIN(N__39198),
            .DOUT(N__39197),
            .PACKAGEPIN(SCK));
    defparam SCK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam SCK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO SCK_ibuf_preio (
            .PADOEN(N__39199),
            .PADOUT(N__39198),
            .PADIN(N__39197),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SCK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ch3_A_ibuf_iopad.PULLUP=1'b1;
    IO_PAD ch3_A_ibuf_iopad (
            .OE(N__39190),
            .DIN(N__39189),
            .DOUT(N__39188),
            .PACKAGEPIN(ch3_A));
    defparam ch3_A_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ch3_A_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ch3_A_ibuf_preio (
            .PADOEN(N__39190),
            .PADOUT(N__39189),
            .PADIN(N__39188),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ch3_A_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ch1_B_ibuf_iopad.PULLUP=1'b1;
    IO_PAD ch1_B_ibuf_iopad (
            .OE(N__39181),
            .DIN(N__39180),
            .DOUT(N__39179),
            .PACKAGEPIN(ch1_B));
    defparam ch1_B_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ch1_B_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ch1_B_ibuf_preio (
            .PADOEN(N__39181),
            .PADOUT(N__39180),
            .PADIN(N__39179),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ch1_B_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PWM2_obuf_iopad (
            .OE(N__39172),
            .DIN(N__39171),
            .DOUT(N__39170),
            .PACKAGEPIN(PWM2));
    defparam PWM2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PWM2_obuf_preio.PIN_TYPE=6'b101001;
    PRE_IO PWM2_obuf_preio (
            .PADOEN(N__39172),
            .PADOUT(N__39171),
            .PADIN(N__39170),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__35463),
            .DIN0(),
            .DOUT0(N__32151),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD MOSI_ibuf_iopad (
            .OE(N__39163),
            .DIN(N__39162),
            .DOUT(N__39161),
            .PACKAGEPIN(MOSI));
    defparam MOSI_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam MOSI_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO MOSI_ibuf_preio (
            .PADOEN(N__39163),
            .PADOUT(N__39162),
            .PADIN(N__39161),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(MOSI_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ch7_B_ibuf_iopad.PULLUP=1'b1;
    IO_PAD ch7_B_ibuf_iopad (
            .OE(N__39154),
            .DIN(N__39153),
            .DOUT(N__39152),
            .PACKAGEPIN(ch7_B));
    defparam ch7_B_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ch7_B_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ch7_B_ibuf_preio (
            .PADOEN(N__39154),
            .PADOUT(N__39153),
            .PADIN(N__39152),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ch7_B_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ch0_A_ibuf_iopad.PULLUP=1'b1;
    IO_PAD ch0_A_ibuf_iopad (
            .OE(N__39145),
            .DIN(N__39144),
            .DOUT(N__39143),
            .PACKAGEPIN(ch0_A));
    defparam ch0_A_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ch0_A_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ch0_A_ibuf_preio (
            .PADOEN(N__39145),
            .PADOUT(N__39144),
            .PADIN(N__39143),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ch0_A_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PWM0_obuf_iopad (
            .OE(N__39136),
            .DIN(N__39135),
            .DOUT(N__39134),
            .PACKAGEPIN(PWM0));
    defparam PWM0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PWM0_obuf_preio.PIN_TYPE=6'b101001;
    PRE_IO PWM0_obuf_preio (
            .PADOEN(N__39136),
            .PADOUT(N__39135),
            .PADIN(N__39134),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__17409),
            .DIN0(),
            .DOUT0(N__17250),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SSEL_ibuf_iopad (
            .OE(N__39127),
            .DIN(N__39126),
            .DOUT(N__39125),
            .PACKAGEPIN(SSEL));
    defparam SSEL_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam SSEL_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO SSEL_ibuf_preio (
            .PADOEN(N__39127),
            .PADOUT(N__39126),
            .PADIN(N__39125),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SSEL_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ch1_A_ibuf_iopad.PULLUP=1'b1;
    IO_PAD ch1_A_ibuf_iopad (
            .OE(N__39118),
            .DIN(N__39117),
            .DOUT(N__39116),
            .PACKAGEPIN(ch1_A));
    defparam ch1_A_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ch1_A_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ch1_A_ibuf_preio (
            .PADOEN(N__39118),
            .PADOUT(N__39117),
            .PADIN(N__39116),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ch1_A_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ch2_A_ibuf_iopad.PULLUP=1'b1;
    IO_PAD ch2_A_ibuf_iopad (
            .OE(N__39109),
            .DIN(N__39108),
            .DOUT(N__39107),
            .PACKAGEPIN(ch2_A));
    defparam ch2_A_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam ch2_A_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO ch2_A_ibuf_preio (
            .PADOEN(N__39109),
            .PADOUT(N__39108),
            .PADIN(N__39107),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(ch2_A_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__9448 (
            .O(N__39090),
            .I(N__39087));
    InMux I__9447 (
            .O(N__39087),
            .I(N__39084));
    LocalMux I__9446 (
            .O(N__39084),
            .I(bit_count_RNIU615_0Z0Z_4));
    CascadeMux I__9445 (
            .O(N__39081),
            .I(bit_count_RNIU615_0Z0Z_4_cascade_));
    InMux I__9444 (
            .O(N__39078),
            .I(N__39075));
    LocalMux I__9443 (
            .O(N__39075),
            .I(N__39072));
    Span4Mux_h I__9442 (
            .O(N__39072),
            .I(N__39069));
    Odrv4 I__9441 (
            .O(N__39069),
            .I(SSELr_RNIGO0FZ0Z_1));
    InMux I__9440 (
            .O(N__39066),
            .I(N__39057));
    InMux I__9439 (
            .O(N__39065),
            .I(N__39057));
    InMux I__9438 (
            .O(N__39064),
            .I(N__39057));
    LocalMux I__9437 (
            .O(N__39057),
            .I(N__39050));
    InMux I__9436 (
            .O(N__39056),
            .I(N__39037));
    InMux I__9435 (
            .O(N__39055),
            .I(N__39037));
    InMux I__9434 (
            .O(N__39054),
            .I(N__39037));
    InMux I__9433 (
            .O(N__39053),
            .I(N__39037));
    Span4Mux_h I__9432 (
            .O(N__39050),
            .I(N__39031));
    InMux I__9431 (
            .O(N__39049),
            .I(N__39024));
    InMux I__9430 (
            .O(N__39048),
            .I(N__39024));
    InMux I__9429 (
            .O(N__39047),
            .I(N__39024));
    InMux I__9428 (
            .O(N__39046),
            .I(N__39021));
    LocalMux I__9427 (
            .O(N__39037),
            .I(N__39018));
    InMux I__9426 (
            .O(N__39036),
            .I(N__39011));
    InMux I__9425 (
            .O(N__39035),
            .I(N__39011));
    InMux I__9424 (
            .O(N__39034),
            .I(N__39011));
    Span4Mux_h I__9423 (
            .O(N__39031),
            .I(N__39006));
    LocalMux I__9422 (
            .O(N__39024),
            .I(N__39006));
    LocalMux I__9421 (
            .O(N__39021),
            .I(SSELrZ0Z_1));
    Odrv12 I__9420 (
            .O(N__39018),
            .I(SSELrZ0Z_1));
    LocalMux I__9419 (
            .O(N__39011),
            .I(SSELrZ0Z_1));
    Odrv4 I__9418 (
            .O(N__39006),
            .I(SSELrZ0Z_1));
    CascadeMux I__9417 (
            .O(N__38997),
            .I(N__38994));
    InMux I__9416 (
            .O(N__38994),
            .I(N__38988));
    InMux I__9415 (
            .O(N__38993),
            .I(N__38988));
    LocalMux I__9414 (
            .O(N__38988),
            .I(un1_bit_count_1_c3));
    InMux I__9413 (
            .O(N__38985),
            .I(N__38979));
    InMux I__9412 (
            .O(N__38984),
            .I(N__38972));
    InMux I__9411 (
            .O(N__38983),
            .I(N__38972));
    InMux I__9410 (
            .O(N__38982),
            .I(N__38972));
    LocalMux I__9409 (
            .O(N__38979),
            .I(bit_countZ0Z_3));
    LocalMux I__9408 (
            .O(N__38972),
            .I(bit_countZ0Z_3));
    InMux I__9407 (
            .O(N__38967),
            .I(N__38962));
    InMux I__9406 (
            .O(N__38966),
            .I(N__38957));
    InMux I__9405 (
            .O(N__38965),
            .I(N__38957));
    LocalMux I__9404 (
            .O(N__38962),
            .I(bit_countZ0Z_4));
    LocalMux I__9403 (
            .O(N__38957),
            .I(bit_countZ0Z_4));
    CascadeMux I__9402 (
            .O(N__38952),
            .I(N__38948));
    InMux I__9401 (
            .O(N__38951),
            .I(N__38943));
    InMux I__9400 (
            .O(N__38948),
            .I(N__38938));
    InMux I__9399 (
            .O(N__38947),
            .I(N__38938));
    InMux I__9398 (
            .O(N__38946),
            .I(N__38934));
    LocalMux I__9397 (
            .O(N__38943),
            .I(N__38929));
    LocalMux I__9396 (
            .O(N__38938),
            .I(N__38926));
    InMux I__9395 (
            .O(N__38937),
            .I(N__38923));
    LocalMux I__9394 (
            .O(N__38934),
            .I(N__38920));
    InMux I__9393 (
            .O(N__38933),
            .I(N__38917));
    InMux I__9392 (
            .O(N__38932),
            .I(N__38914));
    Span4Mux_v I__9391 (
            .O(N__38929),
            .I(N__38905));
    Span4Mux_v I__9390 (
            .O(N__38926),
            .I(N__38905));
    LocalMux I__9389 (
            .O(N__38923),
            .I(N__38902));
    Span4Mux_h I__9388 (
            .O(N__38920),
            .I(N__38893));
    LocalMux I__9387 (
            .O(N__38917),
            .I(N__38893));
    LocalMux I__9386 (
            .O(N__38914),
            .I(N__38893));
    InMux I__9385 (
            .O(N__38913),
            .I(N__38890));
    InMux I__9384 (
            .O(N__38912),
            .I(N__38887));
    CascadeMux I__9383 (
            .O(N__38911),
            .I(N__38884));
    CascadeMux I__9382 (
            .O(N__38910),
            .I(N__38880));
    Span4Mux_h I__9381 (
            .O(N__38905),
            .I(N__38872));
    Span4Mux_h I__9380 (
            .O(N__38902),
            .I(N__38872));
    InMux I__9379 (
            .O(N__38901),
            .I(N__38869));
    InMux I__9378 (
            .O(N__38900),
            .I(N__38866));
    Span4Mux_v I__9377 (
            .O(N__38893),
            .I(N__38857));
    LocalMux I__9376 (
            .O(N__38890),
            .I(N__38857));
    LocalMux I__9375 (
            .O(N__38887),
            .I(N__38857));
    InMux I__9374 (
            .O(N__38884),
            .I(N__38852));
    InMux I__9373 (
            .O(N__38883),
            .I(N__38852));
    InMux I__9372 (
            .O(N__38880),
            .I(N__38847));
    InMux I__9371 (
            .O(N__38879),
            .I(N__38847));
    InMux I__9370 (
            .O(N__38878),
            .I(N__38842));
    InMux I__9369 (
            .O(N__38877),
            .I(N__38842));
    Span4Mux_h I__9368 (
            .O(N__38872),
            .I(N__38837));
    LocalMux I__9367 (
            .O(N__38869),
            .I(N__38837));
    LocalMux I__9366 (
            .O(N__38866),
            .I(N__38834));
    InMux I__9365 (
            .O(N__38865),
            .I(N__38831));
    InMux I__9364 (
            .O(N__38864),
            .I(N__38828));
    Span4Mux_h I__9363 (
            .O(N__38857),
            .I(N__38825));
    LocalMux I__9362 (
            .O(N__38852),
            .I(N__38818));
    LocalMux I__9361 (
            .O(N__38847),
            .I(N__38818));
    LocalMux I__9360 (
            .O(N__38842),
            .I(N__38818));
    Odrv4 I__9359 (
            .O(N__38837),
            .I(un1_OutReg51_4_0_i_o3_3));
    Odrv4 I__9358 (
            .O(N__38834),
            .I(un1_OutReg51_4_0_i_o3_3));
    LocalMux I__9357 (
            .O(N__38831),
            .I(un1_OutReg51_4_0_i_o3_3));
    LocalMux I__9356 (
            .O(N__38828),
            .I(un1_OutReg51_4_0_i_o3_3));
    Odrv4 I__9355 (
            .O(N__38825),
            .I(un1_OutReg51_4_0_i_o3_3));
    Odrv12 I__9354 (
            .O(N__38818),
            .I(un1_OutReg51_4_0_i_o3_3));
    CascadeMux I__9353 (
            .O(N__38805),
            .I(N__38802));
    InMux I__9352 (
            .O(N__38802),
            .I(N__38799));
    LocalMux I__9351 (
            .O(N__38799),
            .I(N__38790));
    InMux I__9350 (
            .O(N__38798),
            .I(N__38787));
    InMux I__9349 (
            .O(N__38797),
            .I(N__38782));
    InMux I__9348 (
            .O(N__38796),
            .I(N__38782));
    InMux I__9347 (
            .O(N__38795),
            .I(N__38777));
    InMux I__9346 (
            .O(N__38794),
            .I(N__38777));
    InMux I__9345 (
            .O(N__38793),
            .I(N__38774));
    Odrv4 I__9344 (
            .O(N__38790),
            .I(SCKrZ0Z_1));
    LocalMux I__9343 (
            .O(N__38787),
            .I(SCKrZ0Z_1));
    LocalMux I__9342 (
            .O(N__38782),
            .I(SCKrZ0Z_1));
    LocalMux I__9341 (
            .O(N__38777),
            .I(SCKrZ0Z_1));
    LocalMux I__9340 (
            .O(N__38774),
            .I(SCKrZ0Z_1));
    CascadeMux I__9339 (
            .O(N__38763),
            .I(N__38755));
    CascadeMux I__9338 (
            .O(N__38762),
            .I(N__38752));
    InMux I__9337 (
            .O(N__38761),
            .I(N__38747));
    InMux I__9336 (
            .O(N__38760),
            .I(N__38747));
    InMux I__9335 (
            .O(N__38759),
            .I(N__38744));
    InMux I__9334 (
            .O(N__38758),
            .I(N__38741));
    InMux I__9333 (
            .O(N__38755),
            .I(N__38738));
    InMux I__9332 (
            .O(N__38752),
            .I(N__38735));
    LocalMux I__9331 (
            .O(N__38747),
            .I(SCKrZ0Z_2));
    LocalMux I__9330 (
            .O(N__38744),
            .I(SCKrZ0Z_2));
    LocalMux I__9329 (
            .O(N__38741),
            .I(SCKrZ0Z_2));
    LocalMux I__9328 (
            .O(N__38738),
            .I(SCKrZ0Z_2));
    LocalMux I__9327 (
            .O(N__38735),
            .I(SCKrZ0Z_2));
    ClkMux I__9326 (
            .O(N__38724),
            .I(N__38172));
    ClkMux I__9325 (
            .O(N__38723),
            .I(N__38172));
    ClkMux I__9324 (
            .O(N__38722),
            .I(N__38172));
    ClkMux I__9323 (
            .O(N__38721),
            .I(N__38172));
    ClkMux I__9322 (
            .O(N__38720),
            .I(N__38172));
    ClkMux I__9321 (
            .O(N__38719),
            .I(N__38172));
    ClkMux I__9320 (
            .O(N__38718),
            .I(N__38172));
    ClkMux I__9319 (
            .O(N__38717),
            .I(N__38172));
    ClkMux I__9318 (
            .O(N__38716),
            .I(N__38172));
    ClkMux I__9317 (
            .O(N__38715),
            .I(N__38172));
    ClkMux I__9316 (
            .O(N__38714),
            .I(N__38172));
    ClkMux I__9315 (
            .O(N__38713),
            .I(N__38172));
    ClkMux I__9314 (
            .O(N__38712),
            .I(N__38172));
    ClkMux I__9313 (
            .O(N__38711),
            .I(N__38172));
    ClkMux I__9312 (
            .O(N__38710),
            .I(N__38172));
    ClkMux I__9311 (
            .O(N__38709),
            .I(N__38172));
    ClkMux I__9310 (
            .O(N__38708),
            .I(N__38172));
    ClkMux I__9309 (
            .O(N__38707),
            .I(N__38172));
    ClkMux I__9308 (
            .O(N__38706),
            .I(N__38172));
    ClkMux I__9307 (
            .O(N__38705),
            .I(N__38172));
    ClkMux I__9306 (
            .O(N__38704),
            .I(N__38172));
    ClkMux I__9305 (
            .O(N__38703),
            .I(N__38172));
    ClkMux I__9304 (
            .O(N__38702),
            .I(N__38172));
    ClkMux I__9303 (
            .O(N__38701),
            .I(N__38172));
    ClkMux I__9302 (
            .O(N__38700),
            .I(N__38172));
    ClkMux I__9301 (
            .O(N__38699),
            .I(N__38172));
    ClkMux I__9300 (
            .O(N__38698),
            .I(N__38172));
    ClkMux I__9299 (
            .O(N__38697),
            .I(N__38172));
    ClkMux I__9298 (
            .O(N__38696),
            .I(N__38172));
    ClkMux I__9297 (
            .O(N__38695),
            .I(N__38172));
    ClkMux I__9296 (
            .O(N__38694),
            .I(N__38172));
    ClkMux I__9295 (
            .O(N__38693),
            .I(N__38172));
    ClkMux I__9294 (
            .O(N__38692),
            .I(N__38172));
    ClkMux I__9293 (
            .O(N__38691),
            .I(N__38172));
    ClkMux I__9292 (
            .O(N__38690),
            .I(N__38172));
    ClkMux I__9291 (
            .O(N__38689),
            .I(N__38172));
    ClkMux I__9290 (
            .O(N__38688),
            .I(N__38172));
    ClkMux I__9289 (
            .O(N__38687),
            .I(N__38172));
    ClkMux I__9288 (
            .O(N__38686),
            .I(N__38172));
    ClkMux I__9287 (
            .O(N__38685),
            .I(N__38172));
    ClkMux I__9286 (
            .O(N__38684),
            .I(N__38172));
    ClkMux I__9285 (
            .O(N__38683),
            .I(N__38172));
    ClkMux I__9284 (
            .O(N__38682),
            .I(N__38172));
    ClkMux I__9283 (
            .O(N__38681),
            .I(N__38172));
    ClkMux I__9282 (
            .O(N__38680),
            .I(N__38172));
    ClkMux I__9281 (
            .O(N__38679),
            .I(N__38172));
    ClkMux I__9280 (
            .O(N__38678),
            .I(N__38172));
    ClkMux I__9279 (
            .O(N__38677),
            .I(N__38172));
    ClkMux I__9278 (
            .O(N__38676),
            .I(N__38172));
    ClkMux I__9277 (
            .O(N__38675),
            .I(N__38172));
    ClkMux I__9276 (
            .O(N__38674),
            .I(N__38172));
    ClkMux I__9275 (
            .O(N__38673),
            .I(N__38172));
    ClkMux I__9274 (
            .O(N__38672),
            .I(N__38172));
    ClkMux I__9273 (
            .O(N__38671),
            .I(N__38172));
    ClkMux I__9272 (
            .O(N__38670),
            .I(N__38172));
    ClkMux I__9271 (
            .O(N__38669),
            .I(N__38172));
    ClkMux I__9270 (
            .O(N__38668),
            .I(N__38172));
    ClkMux I__9269 (
            .O(N__38667),
            .I(N__38172));
    ClkMux I__9268 (
            .O(N__38666),
            .I(N__38172));
    ClkMux I__9267 (
            .O(N__38665),
            .I(N__38172));
    ClkMux I__9266 (
            .O(N__38664),
            .I(N__38172));
    ClkMux I__9265 (
            .O(N__38663),
            .I(N__38172));
    ClkMux I__9264 (
            .O(N__38662),
            .I(N__38172));
    ClkMux I__9263 (
            .O(N__38661),
            .I(N__38172));
    ClkMux I__9262 (
            .O(N__38660),
            .I(N__38172));
    ClkMux I__9261 (
            .O(N__38659),
            .I(N__38172));
    ClkMux I__9260 (
            .O(N__38658),
            .I(N__38172));
    ClkMux I__9259 (
            .O(N__38657),
            .I(N__38172));
    ClkMux I__9258 (
            .O(N__38656),
            .I(N__38172));
    ClkMux I__9257 (
            .O(N__38655),
            .I(N__38172));
    ClkMux I__9256 (
            .O(N__38654),
            .I(N__38172));
    ClkMux I__9255 (
            .O(N__38653),
            .I(N__38172));
    ClkMux I__9254 (
            .O(N__38652),
            .I(N__38172));
    ClkMux I__9253 (
            .O(N__38651),
            .I(N__38172));
    ClkMux I__9252 (
            .O(N__38650),
            .I(N__38172));
    ClkMux I__9251 (
            .O(N__38649),
            .I(N__38172));
    ClkMux I__9250 (
            .O(N__38648),
            .I(N__38172));
    ClkMux I__9249 (
            .O(N__38647),
            .I(N__38172));
    ClkMux I__9248 (
            .O(N__38646),
            .I(N__38172));
    ClkMux I__9247 (
            .O(N__38645),
            .I(N__38172));
    ClkMux I__9246 (
            .O(N__38644),
            .I(N__38172));
    ClkMux I__9245 (
            .O(N__38643),
            .I(N__38172));
    ClkMux I__9244 (
            .O(N__38642),
            .I(N__38172));
    ClkMux I__9243 (
            .O(N__38641),
            .I(N__38172));
    ClkMux I__9242 (
            .O(N__38640),
            .I(N__38172));
    ClkMux I__9241 (
            .O(N__38639),
            .I(N__38172));
    ClkMux I__9240 (
            .O(N__38638),
            .I(N__38172));
    ClkMux I__9239 (
            .O(N__38637),
            .I(N__38172));
    ClkMux I__9238 (
            .O(N__38636),
            .I(N__38172));
    ClkMux I__9237 (
            .O(N__38635),
            .I(N__38172));
    ClkMux I__9236 (
            .O(N__38634),
            .I(N__38172));
    ClkMux I__9235 (
            .O(N__38633),
            .I(N__38172));
    ClkMux I__9234 (
            .O(N__38632),
            .I(N__38172));
    ClkMux I__9233 (
            .O(N__38631),
            .I(N__38172));
    ClkMux I__9232 (
            .O(N__38630),
            .I(N__38172));
    ClkMux I__9231 (
            .O(N__38629),
            .I(N__38172));
    ClkMux I__9230 (
            .O(N__38628),
            .I(N__38172));
    ClkMux I__9229 (
            .O(N__38627),
            .I(N__38172));
    ClkMux I__9228 (
            .O(N__38626),
            .I(N__38172));
    ClkMux I__9227 (
            .O(N__38625),
            .I(N__38172));
    ClkMux I__9226 (
            .O(N__38624),
            .I(N__38172));
    ClkMux I__9225 (
            .O(N__38623),
            .I(N__38172));
    ClkMux I__9224 (
            .O(N__38622),
            .I(N__38172));
    ClkMux I__9223 (
            .O(N__38621),
            .I(N__38172));
    ClkMux I__9222 (
            .O(N__38620),
            .I(N__38172));
    ClkMux I__9221 (
            .O(N__38619),
            .I(N__38172));
    ClkMux I__9220 (
            .O(N__38618),
            .I(N__38172));
    ClkMux I__9219 (
            .O(N__38617),
            .I(N__38172));
    ClkMux I__9218 (
            .O(N__38616),
            .I(N__38172));
    ClkMux I__9217 (
            .O(N__38615),
            .I(N__38172));
    ClkMux I__9216 (
            .O(N__38614),
            .I(N__38172));
    ClkMux I__9215 (
            .O(N__38613),
            .I(N__38172));
    ClkMux I__9214 (
            .O(N__38612),
            .I(N__38172));
    ClkMux I__9213 (
            .O(N__38611),
            .I(N__38172));
    ClkMux I__9212 (
            .O(N__38610),
            .I(N__38172));
    ClkMux I__9211 (
            .O(N__38609),
            .I(N__38172));
    ClkMux I__9210 (
            .O(N__38608),
            .I(N__38172));
    ClkMux I__9209 (
            .O(N__38607),
            .I(N__38172));
    ClkMux I__9208 (
            .O(N__38606),
            .I(N__38172));
    ClkMux I__9207 (
            .O(N__38605),
            .I(N__38172));
    ClkMux I__9206 (
            .O(N__38604),
            .I(N__38172));
    ClkMux I__9205 (
            .O(N__38603),
            .I(N__38172));
    ClkMux I__9204 (
            .O(N__38602),
            .I(N__38172));
    ClkMux I__9203 (
            .O(N__38601),
            .I(N__38172));
    ClkMux I__9202 (
            .O(N__38600),
            .I(N__38172));
    ClkMux I__9201 (
            .O(N__38599),
            .I(N__38172));
    ClkMux I__9200 (
            .O(N__38598),
            .I(N__38172));
    ClkMux I__9199 (
            .O(N__38597),
            .I(N__38172));
    ClkMux I__9198 (
            .O(N__38596),
            .I(N__38172));
    ClkMux I__9197 (
            .O(N__38595),
            .I(N__38172));
    ClkMux I__9196 (
            .O(N__38594),
            .I(N__38172));
    ClkMux I__9195 (
            .O(N__38593),
            .I(N__38172));
    ClkMux I__9194 (
            .O(N__38592),
            .I(N__38172));
    ClkMux I__9193 (
            .O(N__38591),
            .I(N__38172));
    ClkMux I__9192 (
            .O(N__38590),
            .I(N__38172));
    ClkMux I__9191 (
            .O(N__38589),
            .I(N__38172));
    ClkMux I__9190 (
            .O(N__38588),
            .I(N__38172));
    ClkMux I__9189 (
            .O(N__38587),
            .I(N__38172));
    ClkMux I__9188 (
            .O(N__38586),
            .I(N__38172));
    ClkMux I__9187 (
            .O(N__38585),
            .I(N__38172));
    ClkMux I__9186 (
            .O(N__38584),
            .I(N__38172));
    ClkMux I__9185 (
            .O(N__38583),
            .I(N__38172));
    ClkMux I__9184 (
            .O(N__38582),
            .I(N__38172));
    ClkMux I__9183 (
            .O(N__38581),
            .I(N__38172));
    ClkMux I__9182 (
            .O(N__38580),
            .I(N__38172));
    ClkMux I__9181 (
            .O(N__38579),
            .I(N__38172));
    ClkMux I__9180 (
            .O(N__38578),
            .I(N__38172));
    ClkMux I__9179 (
            .O(N__38577),
            .I(N__38172));
    ClkMux I__9178 (
            .O(N__38576),
            .I(N__38172));
    ClkMux I__9177 (
            .O(N__38575),
            .I(N__38172));
    ClkMux I__9176 (
            .O(N__38574),
            .I(N__38172));
    ClkMux I__9175 (
            .O(N__38573),
            .I(N__38172));
    ClkMux I__9174 (
            .O(N__38572),
            .I(N__38172));
    ClkMux I__9173 (
            .O(N__38571),
            .I(N__38172));
    ClkMux I__9172 (
            .O(N__38570),
            .I(N__38172));
    ClkMux I__9171 (
            .O(N__38569),
            .I(N__38172));
    ClkMux I__9170 (
            .O(N__38568),
            .I(N__38172));
    ClkMux I__9169 (
            .O(N__38567),
            .I(N__38172));
    ClkMux I__9168 (
            .O(N__38566),
            .I(N__38172));
    ClkMux I__9167 (
            .O(N__38565),
            .I(N__38172));
    ClkMux I__9166 (
            .O(N__38564),
            .I(N__38172));
    ClkMux I__9165 (
            .O(N__38563),
            .I(N__38172));
    ClkMux I__9164 (
            .O(N__38562),
            .I(N__38172));
    ClkMux I__9163 (
            .O(N__38561),
            .I(N__38172));
    ClkMux I__9162 (
            .O(N__38560),
            .I(N__38172));
    ClkMux I__9161 (
            .O(N__38559),
            .I(N__38172));
    ClkMux I__9160 (
            .O(N__38558),
            .I(N__38172));
    ClkMux I__9159 (
            .O(N__38557),
            .I(N__38172));
    ClkMux I__9158 (
            .O(N__38556),
            .I(N__38172));
    ClkMux I__9157 (
            .O(N__38555),
            .I(N__38172));
    ClkMux I__9156 (
            .O(N__38554),
            .I(N__38172));
    ClkMux I__9155 (
            .O(N__38553),
            .I(N__38172));
    ClkMux I__9154 (
            .O(N__38552),
            .I(N__38172));
    ClkMux I__9153 (
            .O(N__38551),
            .I(N__38172));
    ClkMux I__9152 (
            .O(N__38550),
            .I(N__38172));
    ClkMux I__9151 (
            .O(N__38549),
            .I(N__38172));
    ClkMux I__9150 (
            .O(N__38548),
            .I(N__38172));
    ClkMux I__9149 (
            .O(N__38547),
            .I(N__38172));
    ClkMux I__9148 (
            .O(N__38546),
            .I(N__38172));
    ClkMux I__9147 (
            .O(N__38545),
            .I(N__38172));
    ClkMux I__9146 (
            .O(N__38544),
            .I(N__38172));
    ClkMux I__9145 (
            .O(N__38543),
            .I(N__38172));
    ClkMux I__9144 (
            .O(N__38542),
            .I(N__38172));
    ClkMux I__9143 (
            .O(N__38541),
            .I(N__38172));
    GlobalMux I__9142 (
            .O(N__38172),
            .I(N__38169));
    gio2CtrlBuf I__9141 (
            .O(N__38169),
            .I(myclk));
    CascadeMux I__9140 (
            .O(N__38166),
            .I(N__38163));
    InMux I__9139 (
            .O(N__38163),
            .I(N__38160));
    LocalMux I__9138 (
            .O(N__38160),
            .I(N__38149));
    InMux I__9137 (
            .O(N__38159),
            .I(N__38146));
    InMux I__9136 (
            .O(N__38158),
            .I(N__38143));
    InMux I__9135 (
            .O(N__38157),
            .I(N__38140));
    InMux I__9134 (
            .O(N__38156),
            .I(N__38132));
    InMux I__9133 (
            .O(N__38155),
            .I(N__38132));
    InMux I__9132 (
            .O(N__38154),
            .I(N__38129));
    InMux I__9131 (
            .O(N__38153),
            .I(N__38126));
    InMux I__9130 (
            .O(N__38152),
            .I(N__38123));
    Span4Mux_h I__9129 (
            .O(N__38149),
            .I(N__38118));
    LocalMux I__9128 (
            .O(N__38146),
            .I(N__38118));
    LocalMux I__9127 (
            .O(N__38143),
            .I(N__38115));
    LocalMux I__9126 (
            .O(N__38140),
            .I(N__38110));
    InMux I__9125 (
            .O(N__38139),
            .I(N__38107));
    InMux I__9124 (
            .O(N__38138),
            .I(N__38104));
    CascadeMux I__9123 (
            .O(N__38137),
            .I(N__38101));
    LocalMux I__9122 (
            .O(N__38132),
            .I(N__38097));
    LocalMux I__9121 (
            .O(N__38129),
            .I(N__38091));
    LocalMux I__9120 (
            .O(N__38126),
            .I(N__38088));
    LocalMux I__9119 (
            .O(N__38123),
            .I(N__38085));
    Span4Mux_v I__9118 (
            .O(N__38118),
            .I(N__38080));
    Span4Mux_h I__9117 (
            .O(N__38115),
            .I(N__38080));
    InMux I__9116 (
            .O(N__38114),
            .I(N__38077));
    InMux I__9115 (
            .O(N__38113),
            .I(N__38074));
    Span4Mux_v I__9114 (
            .O(N__38110),
            .I(N__38067));
    LocalMux I__9113 (
            .O(N__38107),
            .I(N__38067));
    LocalMux I__9112 (
            .O(N__38104),
            .I(N__38067));
    InMux I__9111 (
            .O(N__38101),
            .I(N__38064));
    InMux I__9110 (
            .O(N__38100),
            .I(N__38061));
    Span4Mux_h I__9109 (
            .O(N__38097),
            .I(N__38058));
    InMux I__9108 (
            .O(N__38096),
            .I(N__38055));
    InMux I__9107 (
            .O(N__38095),
            .I(N__38052));
    InMux I__9106 (
            .O(N__38094),
            .I(N__38049));
    Span4Mux_h I__9105 (
            .O(N__38091),
            .I(N__38042));
    Span4Mux_h I__9104 (
            .O(N__38088),
            .I(N__38042));
    Span4Mux_h I__9103 (
            .O(N__38085),
            .I(N__38042));
    Span4Mux_h I__9102 (
            .O(N__38080),
            .I(N__38037));
    LocalMux I__9101 (
            .O(N__38077),
            .I(N__38037));
    LocalMux I__9100 (
            .O(N__38074),
            .I(N__38030));
    Span4Mux_h I__9099 (
            .O(N__38067),
            .I(N__38030));
    LocalMux I__9098 (
            .O(N__38064),
            .I(N__38030));
    LocalMux I__9097 (
            .O(N__38061),
            .I(data_receivedZ0Z_0));
    Odrv4 I__9096 (
            .O(N__38058),
            .I(data_receivedZ0Z_0));
    LocalMux I__9095 (
            .O(N__38055),
            .I(data_receivedZ0Z_0));
    LocalMux I__9094 (
            .O(N__38052),
            .I(data_receivedZ0Z_0));
    LocalMux I__9093 (
            .O(N__38049),
            .I(data_receivedZ0Z_0));
    Odrv4 I__9092 (
            .O(N__38042),
            .I(data_receivedZ0Z_0));
    Odrv4 I__9091 (
            .O(N__38037),
            .I(data_receivedZ0Z_0));
    Odrv4 I__9090 (
            .O(N__38030),
            .I(data_receivedZ0Z_0));
    InMux I__9089 (
            .O(N__38013),
            .I(N__38010));
    LocalMux I__9088 (
            .O(N__38010),
            .I(N__38007));
    Span4Mux_v I__9087 (
            .O(N__38007),
            .I(N__38004));
    Odrv4 I__9086 (
            .O(N__38004),
            .I(OutReg_0_5_i_m3_ns_1_8));
    InMux I__9085 (
            .O(N__38001),
            .I(N__37998));
    LocalMux I__9084 (
            .O(N__37998),
            .I(OutReg_esr_RNO_2Z0Z_8));
    InMux I__9083 (
            .O(N__37995),
            .I(N__37992));
    LocalMux I__9082 (
            .O(N__37992),
            .I(N__37989));
    Odrv4 I__9081 (
            .O(N__37989),
            .I(SSELrZ0Z_0));
    InMux I__9080 (
            .O(N__37986),
            .I(N__37977));
    InMux I__9079 (
            .O(N__37985),
            .I(N__37977));
    InMux I__9078 (
            .O(N__37984),
            .I(N__37977));
    LocalMux I__9077 (
            .O(N__37977),
            .I(N__37974));
    Odrv12 I__9076 (
            .O(N__37974),
            .I(SSELrZ0Z_2));
    InMux I__9075 (
            .O(N__37971),
            .I(N__37968));
    LocalMux I__9074 (
            .O(N__37968),
            .I(N__37965));
    Odrv4 I__9073 (
            .O(N__37965),
            .I(SCK_c));
    InMux I__9072 (
            .O(N__37962),
            .I(N__37957));
    InMux I__9071 (
            .O(N__37961),
            .I(N__37954));
    InMux I__9070 (
            .O(N__37960),
            .I(N__37951));
    LocalMux I__9069 (
            .O(N__37957),
            .I(N__37946));
    LocalMux I__9068 (
            .O(N__37954),
            .I(N__37946));
    LocalMux I__9067 (
            .O(N__37951),
            .I(bit_countZ0Z_2));
    Odrv4 I__9066 (
            .O(N__37946),
            .I(bit_countZ0Z_2));
    IoInMux I__9065 (
            .O(N__37941),
            .I(N__37938));
    LocalMux I__9064 (
            .O(N__37938),
            .I(N__37935));
    IoSpan4Mux I__9063 (
            .O(N__37935),
            .I(N__37932));
    Sp12to4 I__9062 (
            .O(N__37932),
            .I(N__37929));
    Odrv12 I__9061 (
            .O(N__37929),
            .I(SCKr_RNIBA7CZ0Z_2));
    CascadeMux I__9060 (
            .O(N__37926),
            .I(SCKr_RNIBA7CZ0Z_2_cascade_));
    IoInMux I__9059 (
            .O(N__37923),
            .I(N__37920));
    LocalMux I__9058 (
            .O(N__37920),
            .I(N__37917));
    Span4Mux_s0_v I__9057 (
            .O(N__37917),
            .I(N__37914));
    Sp12to4 I__9056 (
            .O(N__37914),
            .I(N__37911));
    Span12Mux_h I__9055 (
            .O(N__37911),
            .I(N__37908));
    Odrv12 I__9054 (
            .O(N__37908),
            .I(N_45_0));
    InMux I__9053 (
            .O(N__37905),
            .I(N__37902));
    LocalMux I__9052 (
            .O(N__37902),
            .I(N__37899));
    Odrv12 I__9051 (
            .O(N__37899),
            .I(SCKrZ0Z_0));
    InMux I__9050 (
            .O(N__37896),
            .I(N__37890));
    InMux I__9049 (
            .O(N__37895),
            .I(N__37890));
    LocalMux I__9048 (
            .O(N__37890),
            .I(un1_bit_count_1_c1));
    InMux I__9047 (
            .O(N__37887),
            .I(N__37881));
    InMux I__9046 (
            .O(N__37886),
            .I(N__37878));
    InMux I__9045 (
            .O(N__37885),
            .I(N__37873));
    InMux I__9044 (
            .O(N__37884),
            .I(N__37873));
    LocalMux I__9043 (
            .O(N__37881),
            .I(N__37868));
    LocalMux I__9042 (
            .O(N__37878),
            .I(N__37868));
    LocalMux I__9041 (
            .O(N__37873),
            .I(bit_countZ0Z_1));
    Odrv4 I__9040 (
            .O(N__37868),
            .I(bit_countZ0Z_1));
    InMux I__9039 (
            .O(N__37863),
            .I(N__37860));
    LocalMux I__9038 (
            .O(N__37860),
            .I(N__37857));
    Span4Mux_v I__9037 (
            .O(N__37857),
            .I(N__37854));
    Sp12to4 I__9036 (
            .O(N__37854),
            .I(N__37851));
    Span12Mux_h I__9035 (
            .O(N__37851),
            .I(N__37848));
    Odrv12 I__9034 (
            .O(N__37848),
            .I(SSEL_c));
    CascadeMux I__9033 (
            .O(N__37845),
            .I(un1_bit_count_1_c1_cascade_));
    InMux I__9032 (
            .O(N__37842),
            .I(N__37839));
    LocalMux I__9031 (
            .O(N__37839),
            .I(N__37836));
    Span4Mux_h I__9030 (
            .O(N__37836),
            .I(N__37833));
    Odrv4 I__9029 (
            .O(N__37833),
            .I(OutReg_ess_RNO_1Z0Z_15));
    InMux I__9028 (
            .O(N__37830),
            .I(N__37827));
    LocalMux I__9027 (
            .O(N__37827),
            .I(N__37824));
    Odrv12 I__9026 (
            .O(N__37824),
            .I(OutReg_ess_RNO_2Z0Z_15));
    InMux I__9025 (
            .O(N__37821),
            .I(N__37818));
    LocalMux I__9024 (
            .O(N__37818),
            .I(N__37815));
    Odrv12 I__9023 (
            .O(N__37815),
            .I(OutReg_ess_RNO_0Z0Z_15));
    InMux I__9022 (
            .O(N__37812),
            .I(N__37807));
    InMux I__9021 (
            .O(N__37811),
            .I(N__37802));
    InMux I__9020 (
            .O(N__37810),
            .I(N__37802));
    LocalMux I__9019 (
            .O(N__37807),
            .I(N__37799));
    LocalMux I__9018 (
            .O(N__37802),
            .I(bit_countZ0Z_0));
    Odrv4 I__9017 (
            .O(N__37799),
            .I(bit_countZ0Z_0));
    InMux I__9016 (
            .O(N__37794),
            .I(N__37791));
    LocalMux I__9015 (
            .O(N__37791),
            .I(N__37788));
    Span4Mux_v I__9014 (
            .O(N__37788),
            .I(N__37784));
    InMux I__9013 (
            .O(N__37787),
            .I(N__37780));
    Span4Mux_h I__9012 (
            .O(N__37784),
            .I(N__37777));
    InMux I__9011 (
            .O(N__37783),
            .I(N__37774));
    LocalMux I__9010 (
            .O(N__37780),
            .I(N__37767));
    Span4Mux_h I__9009 (
            .O(N__37777),
            .I(N__37767));
    LocalMux I__9008 (
            .O(N__37774),
            .I(N__37767));
    Odrv4 I__9007 (
            .O(N__37767),
            .I(dataRead6_8));
    InMux I__9006 (
            .O(N__37764),
            .I(N__37756));
    InMux I__9005 (
            .O(N__37763),
            .I(N__37749));
    InMux I__9004 (
            .O(N__37762),
            .I(N__37749));
    InMux I__9003 (
            .O(N__37761),
            .I(N__37749));
    InMux I__9002 (
            .O(N__37760),
            .I(N__37745));
    InMux I__9001 (
            .O(N__37759),
            .I(N__37738));
    LocalMux I__9000 (
            .O(N__37756),
            .I(N__37734));
    LocalMux I__8999 (
            .O(N__37749),
            .I(N__37731));
    InMux I__8998 (
            .O(N__37748),
            .I(N__37728));
    LocalMux I__8997 (
            .O(N__37745),
            .I(N__37725));
    InMux I__8996 (
            .O(N__37744),
            .I(N__37722));
    InMux I__8995 (
            .O(N__37743),
            .I(N__37719));
    InMux I__8994 (
            .O(N__37742),
            .I(N__37716));
    InMux I__8993 (
            .O(N__37741),
            .I(N__37713));
    LocalMux I__8992 (
            .O(N__37738),
            .I(N__37709));
    InMux I__8991 (
            .O(N__37737),
            .I(N__37705));
    Span4Mux_v I__8990 (
            .O(N__37734),
            .I(N__37694));
    Span4Mux_h I__8989 (
            .O(N__37731),
            .I(N__37694));
    LocalMux I__8988 (
            .O(N__37728),
            .I(N__37694));
    Span4Mux_h I__8987 (
            .O(N__37725),
            .I(N__37689));
    LocalMux I__8986 (
            .O(N__37722),
            .I(N__37689));
    LocalMux I__8985 (
            .O(N__37719),
            .I(N__37686));
    LocalMux I__8984 (
            .O(N__37716),
            .I(N__37681));
    LocalMux I__8983 (
            .O(N__37713),
            .I(N__37681));
    InMux I__8982 (
            .O(N__37712),
            .I(N__37678));
    Span4Mux_h I__8981 (
            .O(N__37709),
            .I(N__37675));
    InMux I__8980 (
            .O(N__37708),
            .I(N__37672));
    LocalMux I__8979 (
            .O(N__37705),
            .I(N__37669));
    InMux I__8978 (
            .O(N__37704),
            .I(N__37666));
    InMux I__8977 (
            .O(N__37703),
            .I(N__37663));
    InMux I__8976 (
            .O(N__37702),
            .I(N__37660));
    InMux I__8975 (
            .O(N__37701),
            .I(N__37657));
    Span4Mux_h I__8974 (
            .O(N__37694),
            .I(N__37654));
    Span4Mux_h I__8973 (
            .O(N__37689),
            .I(N__37647));
    Span4Mux_h I__8972 (
            .O(N__37686),
            .I(N__37647));
    Span4Mux_h I__8971 (
            .O(N__37681),
            .I(N__37647));
    LocalMux I__8970 (
            .O(N__37678),
            .I(N__37640));
    Span4Mux_h I__8969 (
            .O(N__37675),
            .I(N__37640));
    LocalMux I__8968 (
            .O(N__37672),
            .I(N__37640));
    Span12Mux_s7_v I__8967 (
            .O(N__37669),
            .I(N__37637));
    LocalMux I__8966 (
            .O(N__37666),
            .I(N__37634));
    LocalMux I__8965 (
            .O(N__37663),
            .I(data_receivedZ0Z_2));
    LocalMux I__8964 (
            .O(N__37660),
            .I(data_receivedZ0Z_2));
    LocalMux I__8963 (
            .O(N__37657),
            .I(data_receivedZ0Z_2));
    Odrv4 I__8962 (
            .O(N__37654),
            .I(data_receivedZ0Z_2));
    Odrv4 I__8961 (
            .O(N__37647),
            .I(data_receivedZ0Z_2));
    Odrv4 I__8960 (
            .O(N__37640),
            .I(data_receivedZ0Z_2));
    Odrv12 I__8959 (
            .O(N__37637),
            .I(data_receivedZ0Z_2));
    Odrv4 I__8958 (
            .O(N__37634),
            .I(data_receivedZ0Z_2));
    CascadeMux I__8957 (
            .O(N__37617),
            .I(N__37614));
    InMux I__8956 (
            .O(N__37614),
            .I(N__37609));
    InMux I__8955 (
            .O(N__37613),
            .I(N__37606));
    InMux I__8954 (
            .O(N__37612),
            .I(N__37603));
    LocalMux I__8953 (
            .O(N__37609),
            .I(N__37600));
    LocalMux I__8952 (
            .O(N__37606),
            .I(N__37595));
    LocalMux I__8951 (
            .O(N__37603),
            .I(N__37595));
    Span4Mux_v I__8950 (
            .O(N__37600),
            .I(N__37592));
    Span4Mux_v I__8949 (
            .O(N__37595),
            .I(N__37589));
    Span4Mux_h I__8948 (
            .O(N__37592),
            .I(N__37586));
    Span4Mux_h I__8947 (
            .O(N__37589),
            .I(N__37583));
    Odrv4 I__8946 (
            .O(N__37586),
            .I(dataRead7_8));
    Odrv4 I__8945 (
            .O(N__37583),
            .I(dataRead7_8));
    InMux I__8944 (
            .O(N__37578),
            .I(N__37575));
    LocalMux I__8943 (
            .O(N__37575),
            .I(N__37572));
    Odrv4 I__8942 (
            .O(N__37572),
            .I(OutReg_0_4_i_m3_ns_1_8));
    InMux I__8941 (
            .O(N__37569),
            .I(N__37566));
    LocalMux I__8940 (
            .O(N__37566),
            .I(N__37553));
    InMux I__8939 (
            .O(N__37565),
            .I(N__37550));
    InMux I__8938 (
            .O(N__37564),
            .I(N__37547));
    InMux I__8937 (
            .O(N__37563),
            .I(N__37544));
    InMux I__8936 (
            .O(N__37562),
            .I(N__37541));
    InMux I__8935 (
            .O(N__37561),
            .I(N__37538));
    InMux I__8934 (
            .O(N__37560),
            .I(N__37534));
    InMux I__8933 (
            .O(N__37559),
            .I(N__37531));
    InMux I__8932 (
            .O(N__37558),
            .I(N__37528));
    InMux I__8931 (
            .O(N__37557),
            .I(N__37525));
    InMux I__8930 (
            .O(N__37556),
            .I(N__37522));
    Span4Mux_h I__8929 (
            .O(N__37553),
            .I(N__37514));
    LocalMux I__8928 (
            .O(N__37550),
            .I(N__37514));
    LocalMux I__8927 (
            .O(N__37547),
            .I(N__37514));
    LocalMux I__8926 (
            .O(N__37544),
            .I(N__37508));
    LocalMux I__8925 (
            .O(N__37541),
            .I(N__37499));
    LocalMux I__8924 (
            .O(N__37538),
            .I(N__37496));
    InMux I__8923 (
            .O(N__37537),
            .I(N__37493));
    LocalMux I__8922 (
            .O(N__37534),
            .I(N__37486));
    LocalMux I__8921 (
            .O(N__37531),
            .I(N__37486));
    LocalMux I__8920 (
            .O(N__37528),
            .I(N__37486));
    LocalMux I__8919 (
            .O(N__37525),
            .I(N__37483));
    LocalMux I__8918 (
            .O(N__37522),
            .I(N__37480));
    InMux I__8917 (
            .O(N__37521),
            .I(N__37477));
    Span4Mux_v I__8916 (
            .O(N__37514),
            .I(N__37474));
    InMux I__8915 (
            .O(N__37513),
            .I(N__37469));
    InMux I__8914 (
            .O(N__37512),
            .I(N__37469));
    InMux I__8913 (
            .O(N__37511),
            .I(N__37466));
    Span12Mux_v I__8912 (
            .O(N__37508),
            .I(N__37463));
    InMux I__8911 (
            .O(N__37507),
            .I(N__37456));
    InMux I__8910 (
            .O(N__37506),
            .I(N__37456));
    InMux I__8909 (
            .O(N__37505),
            .I(N__37456));
    InMux I__8908 (
            .O(N__37504),
            .I(N__37449));
    InMux I__8907 (
            .O(N__37503),
            .I(N__37449));
    InMux I__8906 (
            .O(N__37502),
            .I(N__37449));
    Span4Mux_h I__8905 (
            .O(N__37499),
            .I(N__37444));
    Span4Mux_h I__8904 (
            .O(N__37496),
            .I(N__37444));
    LocalMux I__8903 (
            .O(N__37493),
            .I(N__37439));
    Span4Mux_h I__8902 (
            .O(N__37486),
            .I(N__37439));
    Span4Mux_h I__8901 (
            .O(N__37483),
            .I(N__37434));
    Span4Mux_h I__8900 (
            .O(N__37480),
            .I(N__37434));
    LocalMux I__8899 (
            .O(N__37477),
            .I(N__37427));
    Span4Mux_h I__8898 (
            .O(N__37474),
            .I(N__37427));
    LocalMux I__8897 (
            .O(N__37469),
            .I(N__37427));
    LocalMux I__8896 (
            .O(N__37466),
            .I(data_receivedZ0Z_1));
    Odrv12 I__8895 (
            .O(N__37463),
            .I(data_receivedZ0Z_1));
    LocalMux I__8894 (
            .O(N__37456),
            .I(data_receivedZ0Z_1));
    LocalMux I__8893 (
            .O(N__37449),
            .I(data_receivedZ0Z_1));
    Odrv4 I__8892 (
            .O(N__37444),
            .I(data_receivedZ0Z_1));
    Odrv4 I__8891 (
            .O(N__37439),
            .I(data_receivedZ0Z_1));
    Odrv4 I__8890 (
            .O(N__37434),
            .I(data_receivedZ0Z_1));
    Odrv4 I__8889 (
            .O(N__37427),
            .I(data_receivedZ0Z_1));
    CascadeMux I__8888 (
            .O(N__37410),
            .I(OutReg_esr_RNO_1Z0Z_8_cascade_));
    InMux I__8887 (
            .O(N__37407),
            .I(N__37404));
    LocalMux I__8886 (
            .O(N__37404),
            .I(N__37401));
    Odrv12 I__8885 (
            .O(N__37401),
            .I(OutRegZ0Z_7));
    CascadeMux I__8884 (
            .O(N__37398),
            .I(OutReg_esr_RNO_0Z0Z_8_cascade_));
    InMux I__8883 (
            .O(N__37395),
            .I(N__37389));
    InMux I__8882 (
            .O(N__37394),
            .I(N__37389));
    LocalMux I__8881 (
            .O(N__37389),
            .I(N__37382));
    InMux I__8880 (
            .O(N__37388),
            .I(N__37375));
    InMux I__8879 (
            .O(N__37387),
            .I(N__37371));
    InMux I__8878 (
            .O(N__37386),
            .I(N__37366));
    InMux I__8877 (
            .O(N__37385),
            .I(N__37366));
    Span4Mux_h I__8876 (
            .O(N__37382),
            .I(N__37363));
    InMux I__8875 (
            .O(N__37381),
            .I(N__37360));
    InMux I__8874 (
            .O(N__37380),
            .I(N__37357));
    InMux I__8873 (
            .O(N__37379),
            .I(N__37352));
    InMux I__8872 (
            .O(N__37378),
            .I(N__37352));
    LocalMux I__8871 (
            .O(N__37375),
            .I(N__37348));
    InMux I__8870 (
            .O(N__37374),
            .I(N__37345));
    LocalMux I__8869 (
            .O(N__37371),
            .I(N__37341));
    LocalMux I__8868 (
            .O(N__37366),
            .I(N__37338));
    Span4Mux_h I__8867 (
            .O(N__37363),
            .I(N__37333));
    LocalMux I__8866 (
            .O(N__37360),
            .I(N__37333));
    LocalMux I__8865 (
            .O(N__37357),
            .I(N__37327));
    LocalMux I__8864 (
            .O(N__37352),
            .I(N__37327));
    InMux I__8863 (
            .O(N__37351),
            .I(N__37324));
    Span4Mux_v I__8862 (
            .O(N__37348),
            .I(N__37317));
    LocalMux I__8861 (
            .O(N__37345),
            .I(N__37317));
    InMux I__8860 (
            .O(N__37344),
            .I(N__37314));
    Span4Mux_h I__8859 (
            .O(N__37341),
            .I(N__37307));
    Span4Mux_h I__8858 (
            .O(N__37338),
            .I(N__37307));
    Span4Mux_h I__8857 (
            .O(N__37333),
            .I(N__37304));
    InMux I__8856 (
            .O(N__37332),
            .I(N__37301));
    Span4Mux_v I__8855 (
            .O(N__37327),
            .I(N__37296));
    LocalMux I__8854 (
            .O(N__37324),
            .I(N__37296));
    InMux I__8853 (
            .O(N__37323),
            .I(N__37293));
    InMux I__8852 (
            .O(N__37322),
            .I(N__37290));
    Span4Mux_h I__8851 (
            .O(N__37317),
            .I(N__37285));
    LocalMux I__8850 (
            .O(N__37314),
            .I(N__37285));
    InMux I__8849 (
            .O(N__37313),
            .I(N__37280));
    InMux I__8848 (
            .O(N__37312),
            .I(N__37280));
    Odrv4 I__8847 (
            .O(N__37307),
            .I(un1_OutReg51_4_0_i_o3_2));
    Odrv4 I__8846 (
            .O(N__37304),
            .I(un1_OutReg51_4_0_i_o3_2));
    LocalMux I__8845 (
            .O(N__37301),
            .I(un1_OutReg51_4_0_i_o3_2));
    Odrv4 I__8844 (
            .O(N__37296),
            .I(un1_OutReg51_4_0_i_o3_2));
    LocalMux I__8843 (
            .O(N__37293),
            .I(un1_OutReg51_4_0_i_o3_2));
    LocalMux I__8842 (
            .O(N__37290),
            .I(un1_OutReg51_4_0_i_o3_2));
    Odrv4 I__8841 (
            .O(N__37285),
            .I(un1_OutReg51_4_0_i_o3_2));
    LocalMux I__8840 (
            .O(N__37280),
            .I(un1_OutReg51_4_0_i_o3_2));
    InMux I__8839 (
            .O(N__37263),
            .I(N__37260));
    LocalMux I__8838 (
            .O(N__37260),
            .I(N__37257));
    Sp12to4 I__8837 (
            .O(N__37257),
            .I(N__37254));
    Odrv12 I__8836 (
            .O(N__37254),
            .I(OutRegZ0Z_8));
    CEMux I__8835 (
            .O(N__37251),
            .I(N__37247));
    CEMux I__8834 (
            .O(N__37250),
            .I(N__37237));
    LocalMux I__8833 (
            .O(N__37247),
            .I(N__37234));
    CEMux I__8832 (
            .O(N__37246),
            .I(N__37231));
    CEMux I__8831 (
            .O(N__37245),
            .I(N__37228));
    CEMux I__8830 (
            .O(N__37244),
            .I(N__37225));
    CEMux I__8829 (
            .O(N__37243),
            .I(N__37221));
    CEMux I__8828 (
            .O(N__37242),
            .I(N__37218));
    CEMux I__8827 (
            .O(N__37241),
            .I(N__37215));
    CEMux I__8826 (
            .O(N__37240),
            .I(N__37212));
    LocalMux I__8825 (
            .O(N__37237),
            .I(N__37207));
    Span4Mux_h I__8824 (
            .O(N__37234),
            .I(N__37202));
    LocalMux I__8823 (
            .O(N__37231),
            .I(N__37202));
    LocalMux I__8822 (
            .O(N__37228),
            .I(N__37197));
    LocalMux I__8821 (
            .O(N__37225),
            .I(N__37197));
    CEMux I__8820 (
            .O(N__37224),
            .I(N__37194));
    LocalMux I__8819 (
            .O(N__37221),
            .I(N__37191));
    LocalMux I__8818 (
            .O(N__37218),
            .I(N__37186));
    LocalMux I__8817 (
            .O(N__37215),
            .I(N__37186));
    LocalMux I__8816 (
            .O(N__37212),
            .I(N__37183));
    CEMux I__8815 (
            .O(N__37211),
            .I(N__37180));
    CEMux I__8814 (
            .O(N__37210),
            .I(N__37177));
    Span4Mux_h I__8813 (
            .O(N__37207),
            .I(N__37174));
    Span4Mux_v I__8812 (
            .O(N__37202),
            .I(N__37171));
    Span4Mux_h I__8811 (
            .O(N__37197),
            .I(N__37168));
    LocalMux I__8810 (
            .O(N__37194),
            .I(N__37165));
    Span4Mux_v I__8809 (
            .O(N__37191),
            .I(N__37160));
    Span4Mux_h I__8808 (
            .O(N__37186),
            .I(N__37160));
    Sp12to4 I__8807 (
            .O(N__37183),
            .I(N__37155));
    LocalMux I__8806 (
            .O(N__37180),
            .I(N__37155));
    LocalMux I__8805 (
            .O(N__37177),
            .I(N__37152));
    Odrv4 I__8804 (
            .O(N__37174),
            .I(N_863_0));
    Odrv4 I__8803 (
            .O(N__37171),
            .I(N_863_0));
    Odrv4 I__8802 (
            .O(N__37168),
            .I(N_863_0));
    Odrv4 I__8801 (
            .O(N__37165),
            .I(N_863_0));
    Odrv4 I__8800 (
            .O(N__37160),
            .I(N_863_0));
    Odrv12 I__8799 (
            .O(N__37155),
            .I(N_863_0));
    Odrv12 I__8798 (
            .O(N__37152),
            .I(N_863_0));
    SRMux I__8797 (
            .O(N__37137),
            .I(N__37125));
    SRMux I__8796 (
            .O(N__37136),
            .I(N__37122));
    SRMux I__8795 (
            .O(N__37135),
            .I(N__37119));
    SRMux I__8794 (
            .O(N__37134),
            .I(N__37116));
    SRMux I__8793 (
            .O(N__37133),
            .I(N__37112));
    SRMux I__8792 (
            .O(N__37132),
            .I(N__37109));
    SRMux I__8791 (
            .O(N__37131),
            .I(N__37106));
    SRMux I__8790 (
            .O(N__37130),
            .I(N__37103));
    SRMux I__8789 (
            .O(N__37129),
            .I(N__37100));
    SRMux I__8788 (
            .O(N__37128),
            .I(N__37096));
    LocalMux I__8787 (
            .O(N__37125),
            .I(N__37093));
    LocalMux I__8786 (
            .O(N__37122),
            .I(N__37090));
    LocalMux I__8785 (
            .O(N__37119),
            .I(N__37087));
    LocalMux I__8784 (
            .O(N__37116),
            .I(N__37084));
    SRMux I__8783 (
            .O(N__37115),
            .I(N__37081));
    LocalMux I__8782 (
            .O(N__37112),
            .I(N__37078));
    LocalMux I__8781 (
            .O(N__37109),
            .I(N__37075));
    LocalMux I__8780 (
            .O(N__37106),
            .I(N__37072));
    LocalMux I__8779 (
            .O(N__37103),
            .I(N__37067));
    LocalMux I__8778 (
            .O(N__37100),
            .I(N__37067));
    SRMux I__8777 (
            .O(N__37099),
            .I(N__37064));
    LocalMux I__8776 (
            .O(N__37096),
            .I(N__37061));
    Span4Mux_h I__8775 (
            .O(N__37093),
            .I(N__37055));
    Span4Mux_h I__8774 (
            .O(N__37090),
            .I(N__37055));
    Span4Mux_v I__8773 (
            .O(N__37087),
            .I(N__37050));
    Span4Mux_h I__8772 (
            .O(N__37084),
            .I(N__37050));
    LocalMux I__8771 (
            .O(N__37081),
            .I(N__37047));
    Span4Mux_h I__8770 (
            .O(N__37078),
            .I(N__37038));
    Span4Mux_v I__8769 (
            .O(N__37075),
            .I(N__37038));
    Span4Mux_v I__8768 (
            .O(N__37072),
            .I(N__37038));
    Span4Mux_h I__8767 (
            .O(N__37067),
            .I(N__37038));
    LocalMux I__8766 (
            .O(N__37064),
            .I(N__37033));
    Span4Mux_h I__8765 (
            .O(N__37061),
            .I(N__37033));
    InMux I__8764 (
            .O(N__37060),
            .I(N__37030));
    Odrv4 I__8763 (
            .O(N__37055),
            .I(OutReg_0_sqmuxa));
    Odrv4 I__8762 (
            .O(N__37050),
            .I(OutReg_0_sqmuxa));
    Odrv4 I__8761 (
            .O(N__37047),
            .I(OutReg_0_sqmuxa));
    Odrv4 I__8760 (
            .O(N__37038),
            .I(OutReg_0_sqmuxa));
    Odrv4 I__8759 (
            .O(N__37033),
            .I(OutReg_0_sqmuxa));
    LocalMux I__8758 (
            .O(N__37030),
            .I(OutReg_0_sqmuxa));
    InMux I__8757 (
            .O(N__37017),
            .I(N__37014));
    LocalMux I__8756 (
            .O(N__37014),
            .I(N__37009));
    InMux I__8755 (
            .O(N__37013),
            .I(N__37006));
    InMux I__8754 (
            .O(N__37012),
            .I(N__37003));
    Span4Mux_v I__8753 (
            .O(N__37009),
            .I(N__37000));
    LocalMux I__8752 (
            .O(N__37006),
            .I(N__36995));
    LocalMux I__8751 (
            .O(N__37003),
            .I(N__36995));
    Sp12to4 I__8750 (
            .O(N__37000),
            .I(N__36992));
    Span4Mux_h I__8749 (
            .O(N__36995),
            .I(N__36989));
    Odrv12 I__8748 (
            .O(N__36992),
            .I(dataRead1_8));
    Odrv4 I__8747 (
            .O(N__36989),
            .I(dataRead1_8));
    InMux I__8746 (
            .O(N__36984),
            .I(N__36981));
    LocalMux I__8745 (
            .O(N__36981),
            .I(N__36977));
    InMux I__8744 (
            .O(N__36980),
            .I(N__36974));
    Span4Mux_v I__8743 (
            .O(N__36977),
            .I(N__36970));
    LocalMux I__8742 (
            .O(N__36974),
            .I(N__36967));
    InMux I__8741 (
            .O(N__36973),
            .I(N__36964));
    Span4Mux_h I__8740 (
            .O(N__36970),
            .I(N__36961));
    Span12Mux_h I__8739 (
            .O(N__36967),
            .I(N__36958));
    LocalMux I__8738 (
            .O(N__36964),
            .I(N__36955));
    Odrv4 I__8737 (
            .O(N__36961),
            .I(dataRead5_8));
    Odrv12 I__8736 (
            .O(N__36958),
            .I(dataRead5_8));
    Odrv4 I__8735 (
            .O(N__36955),
            .I(dataRead5_8));
    IoInMux I__8734 (
            .O(N__36948),
            .I(N__36945));
    LocalMux I__8733 (
            .O(N__36945),
            .I(PWM3_obufLegalizeSB_DFFNet));
    IoInMux I__8732 (
            .O(N__36942),
            .I(N__36939));
    LocalMux I__8731 (
            .O(N__36939),
            .I(MISO_obufLegalizeSB_DFFNet));
    ClkMux I__8730 (
            .O(N__36936),
            .I(N__36933));
    LocalMux I__8729 (
            .O(N__36933),
            .I(N__36929));
    ClkMux I__8728 (
            .O(N__36932),
            .I(N__36926));
    Span4Mux_h I__8727 (
            .O(N__36929),
            .I(N__36920));
    LocalMux I__8726 (
            .O(N__36926),
            .I(N__36920));
    ClkMux I__8725 (
            .O(N__36925),
            .I(N__36917));
    Span4Mux_h I__8724 (
            .O(N__36920),
            .I(N__36913));
    LocalMux I__8723 (
            .O(N__36917),
            .I(N__36910));
    ClkMux I__8722 (
            .O(N__36916),
            .I(N__36907));
    Span4Mux_h I__8721 (
            .O(N__36913),
            .I(N__36899));
    Span4Mux_h I__8720 (
            .O(N__36910),
            .I(N__36899));
    LocalMux I__8719 (
            .O(N__36907),
            .I(N__36899));
    ClkMux I__8718 (
            .O(N__36906),
            .I(N__36896));
    Sp12to4 I__8717 (
            .O(N__36899),
            .I(N__36893));
    LocalMux I__8716 (
            .O(N__36896),
            .I(N__36890));
    Span12Mux_h I__8715 (
            .O(N__36893),
            .I(N__36887));
    Span4Mux_h I__8714 (
            .O(N__36890),
            .I(N__36884));
    Span12Mux_v I__8713 (
            .O(N__36887),
            .I(N__36881));
    Span4Mux_h I__8712 (
            .O(N__36884),
            .I(N__36878));
    Odrv12 I__8711 (
            .O(N__36881),
            .I(internalOscilatorOutputNet));
    Odrv4 I__8710 (
            .O(N__36878),
            .I(internalOscilatorOutputNet));
    InMux I__8709 (
            .O(N__36873),
            .I(N__36868));
    InMux I__8708 (
            .O(N__36872),
            .I(N__36865));
    InMux I__8707 (
            .O(N__36871),
            .I(N__36862));
    LocalMux I__8706 (
            .O(N__36868),
            .I(N__36859));
    LocalMux I__8705 (
            .O(N__36865),
            .I(N__36856));
    LocalMux I__8704 (
            .O(N__36862),
            .I(N__36853));
    Span4Mux_v I__8703 (
            .O(N__36859),
            .I(N__36850));
    Span4Mux_h I__8702 (
            .O(N__36856),
            .I(N__36847));
    Span4Mux_h I__8701 (
            .O(N__36853),
            .I(N__36844));
    Span4Mux_h I__8700 (
            .O(N__36850),
            .I(N__36841));
    Sp12to4 I__8699 (
            .O(N__36847),
            .I(N__36838));
    Odrv4 I__8698 (
            .O(N__36844),
            .I(dataRead5_5));
    Odrv4 I__8697 (
            .O(N__36841),
            .I(dataRead5_5));
    Odrv12 I__8696 (
            .O(N__36838),
            .I(dataRead5_5));
    CascadeMux I__8695 (
            .O(N__36831),
            .I(N__36828));
    InMux I__8694 (
            .O(N__36828),
            .I(N__36824));
    InMux I__8693 (
            .O(N__36827),
            .I(N__36821));
    LocalMux I__8692 (
            .O(N__36824),
            .I(N__36818));
    LocalMux I__8691 (
            .O(N__36821),
            .I(N__36814));
    Span4Mux_h I__8690 (
            .O(N__36818),
            .I(N__36811));
    InMux I__8689 (
            .O(N__36817),
            .I(N__36808));
    Span4Mux_v I__8688 (
            .O(N__36814),
            .I(N__36805));
    Span4Mux_h I__8687 (
            .O(N__36811),
            .I(N__36800));
    LocalMux I__8686 (
            .O(N__36808),
            .I(N__36800));
    Odrv4 I__8685 (
            .O(N__36805),
            .I(dataRead1_5));
    Odrv4 I__8684 (
            .O(N__36800),
            .I(dataRead1_5));
    InMux I__8683 (
            .O(N__36795),
            .I(N__36792));
    LocalMux I__8682 (
            .O(N__36792),
            .I(N__36789));
    Span4Mux_v I__8681 (
            .O(N__36789),
            .I(N__36786));
    Odrv4 I__8680 (
            .O(N__36786),
            .I(OutReg_0_5_i_m3_ns_1_5));
    InMux I__8679 (
            .O(N__36783),
            .I(N__36780));
    LocalMux I__8678 (
            .O(N__36780),
            .I(N__36777));
    Span4Mux_v I__8677 (
            .O(N__36777),
            .I(N__36773));
    InMux I__8676 (
            .O(N__36776),
            .I(N__36770));
    Span4Mux_h I__8675 (
            .O(N__36773),
            .I(N__36767));
    LocalMux I__8674 (
            .O(N__36770),
            .I(N__36763));
    Span4Mux_h I__8673 (
            .O(N__36767),
            .I(N__36760));
    InMux I__8672 (
            .O(N__36766),
            .I(N__36757));
    Odrv12 I__8671 (
            .O(N__36763),
            .I(dataRead6_5));
    Odrv4 I__8670 (
            .O(N__36760),
            .I(dataRead6_5));
    LocalMux I__8669 (
            .O(N__36757),
            .I(dataRead6_5));
    CascadeMux I__8668 (
            .O(N__36750),
            .I(N__36747));
    InMux I__8667 (
            .O(N__36747),
            .I(N__36743));
    InMux I__8666 (
            .O(N__36746),
            .I(N__36740));
    LocalMux I__8665 (
            .O(N__36743),
            .I(N__36736));
    LocalMux I__8664 (
            .O(N__36740),
            .I(N__36733));
    InMux I__8663 (
            .O(N__36739),
            .I(N__36730));
    Span4Mux_v I__8662 (
            .O(N__36736),
            .I(N__36727));
    Span4Mux_h I__8661 (
            .O(N__36733),
            .I(N__36722));
    LocalMux I__8660 (
            .O(N__36730),
            .I(N__36722));
    Span4Mux_h I__8659 (
            .O(N__36727),
            .I(N__36719));
    Span4Mux_v I__8658 (
            .O(N__36722),
            .I(N__36716));
    Odrv4 I__8657 (
            .O(N__36719),
            .I(dataRead7_5));
    Odrv4 I__8656 (
            .O(N__36716),
            .I(dataRead7_5));
    InMux I__8655 (
            .O(N__36711),
            .I(N__36708));
    LocalMux I__8654 (
            .O(N__36708),
            .I(N__36705));
    Span4Mux_v I__8653 (
            .O(N__36705),
            .I(N__36702));
    Span4Mux_h I__8652 (
            .O(N__36702),
            .I(N__36699));
    Odrv4 I__8651 (
            .O(N__36699),
            .I(OutReg_0_4_i_m3_ns_1_5));
    CascadeMux I__8650 (
            .O(N__36696),
            .I(OutReg_ess_RNO_1Z0Z_5_cascade_));
    InMux I__8649 (
            .O(N__36693),
            .I(N__36690));
    LocalMux I__8648 (
            .O(N__36690),
            .I(OutReg_ess_RNO_2Z0Z_5));
    InMux I__8647 (
            .O(N__36687),
            .I(N__36684));
    LocalMux I__8646 (
            .O(N__36684),
            .I(OutReg_ess_RNO_0Z0Z_5));
    CascadeMux I__8645 (
            .O(N__36681),
            .I(N__36678));
    InMux I__8644 (
            .O(N__36678),
            .I(N__36675));
    LocalMux I__8643 (
            .O(N__36675),
            .I(N__36672));
    Span4Mux_h I__8642 (
            .O(N__36672),
            .I(N__36669));
    Odrv4 I__8641 (
            .O(N__36669),
            .I(OutRegZ0Z_4));
    InMux I__8640 (
            .O(N__36666),
            .I(N__36663));
    LocalMux I__8639 (
            .O(N__36663),
            .I(N__36660));
    Span4Mux_h I__8638 (
            .O(N__36660),
            .I(N__36657));
    Odrv4 I__8637 (
            .O(N__36657),
            .I(OutRegZ0Z_5));
    InMux I__8636 (
            .O(N__36654),
            .I(N__36651));
    LocalMux I__8635 (
            .O(N__36651),
            .I(N__36648));
    Span4Mux_h I__8634 (
            .O(N__36648),
            .I(N__36645));
    Odrv4 I__8633 (
            .O(N__36645),
            .I(OutRegZ0Z_15));
    CascadeMux I__8632 (
            .O(N__36642),
            .I(dataOut_RNOZ0Z_0_cascade_));
    IoInMux I__8631 (
            .O(N__36639),
            .I(N__36636));
    LocalMux I__8630 (
            .O(N__36636),
            .I(N__36633));
    Span4Mux_s2_v I__8629 (
            .O(N__36633),
            .I(N__36630));
    Span4Mux_v I__8628 (
            .O(N__36630),
            .I(N__36626));
    InMux I__8627 (
            .O(N__36629),
            .I(N__36623));
    Odrv4 I__8626 (
            .O(N__36626),
            .I(MISO_c));
    LocalMux I__8625 (
            .O(N__36623),
            .I(MISO_c));
    InMux I__8624 (
            .O(N__36618),
            .I(N__36613));
    InMux I__8623 (
            .O(N__36617),
            .I(N__36610));
    InMux I__8622 (
            .O(N__36616),
            .I(N__36607));
    LocalMux I__8621 (
            .O(N__36613),
            .I(N__36604));
    LocalMux I__8620 (
            .O(N__36610),
            .I(\PWMInstance2.periodCounterZ0Z_14 ));
    LocalMux I__8619 (
            .O(N__36607),
            .I(\PWMInstance2.periodCounterZ0Z_14 ));
    Odrv4 I__8618 (
            .O(N__36604),
            .I(\PWMInstance2.periodCounterZ0Z_14 ));
    InMux I__8617 (
            .O(N__36597),
            .I(N__36592));
    InMux I__8616 (
            .O(N__36596),
            .I(N__36589));
    InMux I__8615 (
            .O(N__36595),
            .I(N__36586));
    LocalMux I__8614 (
            .O(N__36592),
            .I(N__36581));
    LocalMux I__8613 (
            .O(N__36589),
            .I(N__36581));
    LocalMux I__8612 (
            .O(N__36586),
            .I(\PWMInstance2.periodCounterZ0Z_2 ));
    Odrv4 I__8611 (
            .O(N__36581),
            .I(\PWMInstance2.periodCounterZ0Z_2 ));
    InMux I__8610 (
            .O(N__36576),
            .I(N__36569));
    InMux I__8609 (
            .O(N__36575),
            .I(N__36569));
    InMux I__8608 (
            .O(N__36574),
            .I(N__36566));
    LocalMux I__8607 (
            .O(N__36569),
            .I(N__36563));
    LocalMux I__8606 (
            .O(N__36566),
            .I(\PWMInstance2.periodCounterZ0Z_4 ));
    Odrv4 I__8605 (
            .O(N__36563),
            .I(\PWMInstance2.periodCounterZ0Z_4 ));
    InMux I__8604 (
            .O(N__36558),
            .I(N__36553));
    InMux I__8603 (
            .O(N__36557),
            .I(N__36550));
    InMux I__8602 (
            .O(N__36556),
            .I(N__36547));
    LocalMux I__8601 (
            .O(N__36553),
            .I(N__36544));
    LocalMux I__8600 (
            .O(N__36550),
            .I(\PWMInstance2.periodCounterZ0Z_12 ));
    LocalMux I__8599 (
            .O(N__36547),
            .I(\PWMInstance2.periodCounterZ0Z_12 ));
    Odrv4 I__8598 (
            .O(N__36544),
            .I(\PWMInstance2.periodCounterZ0Z_12 ));
    CascadeMux I__8597 (
            .O(N__36537),
            .I(\PWMInstance2.un1_periodCounter12_1_0_a2_0_0_cascade_ ));
    InMux I__8596 (
            .O(N__36534),
            .I(N__36531));
    LocalMux I__8595 (
            .O(N__36531),
            .I(N__36528));
    Odrv4 I__8594 (
            .O(N__36528),
            .I(\PWMInstance2.un1_periodCounter12_1_0_a2_0_12 ));
    InMux I__8593 (
            .O(N__36525),
            .I(N__36522));
    LocalMux I__8592 (
            .O(N__36522),
            .I(N__36518));
    InMux I__8591 (
            .O(N__36521),
            .I(N__36515));
    Span4Mux_s2_v I__8590 (
            .O(N__36518),
            .I(N__36507));
    LocalMux I__8589 (
            .O(N__36515),
            .I(N__36507));
    InMux I__8588 (
            .O(N__36514),
            .I(N__36504));
    InMux I__8587 (
            .O(N__36513),
            .I(N__36498));
    InMux I__8586 (
            .O(N__36512),
            .I(N__36495));
    Span4Mux_h I__8585 (
            .O(N__36507),
            .I(N__36489));
    LocalMux I__8584 (
            .O(N__36504),
            .I(N__36489));
    InMux I__8583 (
            .O(N__36503),
            .I(N__36480));
    InMux I__8582 (
            .O(N__36502),
            .I(N__36477));
    InMux I__8581 (
            .O(N__36501),
            .I(N__36474));
    LocalMux I__8580 (
            .O(N__36498),
            .I(N__36471));
    LocalMux I__8579 (
            .O(N__36495),
            .I(N__36468));
    InMux I__8578 (
            .O(N__36494),
            .I(N__36465));
    Span4Mux_v I__8577 (
            .O(N__36489),
            .I(N__36462));
    InMux I__8576 (
            .O(N__36488),
            .I(N__36451));
    InMux I__8575 (
            .O(N__36487),
            .I(N__36451));
    InMux I__8574 (
            .O(N__36486),
            .I(N__36451));
    InMux I__8573 (
            .O(N__36485),
            .I(N__36451));
    InMux I__8572 (
            .O(N__36484),
            .I(N__36451));
    CascadeMux I__8571 (
            .O(N__36483),
            .I(N__36448));
    LocalMux I__8570 (
            .O(N__36480),
            .I(N__36445));
    LocalMux I__8569 (
            .O(N__36477),
            .I(N__36442));
    LocalMux I__8568 (
            .O(N__36474),
            .I(N__36439));
    Span4Mux_v I__8567 (
            .O(N__36471),
            .I(N__36435));
    Span4Mux_v I__8566 (
            .O(N__36468),
            .I(N__36430));
    LocalMux I__8565 (
            .O(N__36465),
            .I(N__36430));
    Span4Mux_h I__8564 (
            .O(N__36462),
            .I(N__36427));
    LocalMux I__8563 (
            .O(N__36451),
            .I(N__36424));
    InMux I__8562 (
            .O(N__36448),
            .I(N__36421));
    Span12Mux_h I__8561 (
            .O(N__36445),
            .I(N__36418));
    Span4Mux_v I__8560 (
            .O(N__36442),
            .I(N__36415));
    Span4Mux_v I__8559 (
            .O(N__36439),
            .I(N__36412));
    InMux I__8558 (
            .O(N__36438),
            .I(N__36409));
    Span4Mux_h I__8557 (
            .O(N__36435),
            .I(N__36402));
    Span4Mux_v I__8556 (
            .O(N__36430),
            .I(N__36402));
    Span4Mux_v I__8555 (
            .O(N__36427),
            .I(N__36402));
    Span4Mux_v I__8554 (
            .O(N__36424),
            .I(N__36397));
    LocalMux I__8553 (
            .O(N__36421),
            .I(N__36397));
    Odrv12 I__8552 (
            .O(N__36418),
            .I(dataWriteZ0Z_4));
    Odrv4 I__8551 (
            .O(N__36415),
            .I(dataWriteZ0Z_4));
    Odrv4 I__8550 (
            .O(N__36412),
            .I(dataWriteZ0Z_4));
    LocalMux I__8549 (
            .O(N__36409),
            .I(dataWriteZ0Z_4));
    Odrv4 I__8548 (
            .O(N__36402),
            .I(dataWriteZ0Z_4));
    Odrv4 I__8547 (
            .O(N__36397),
            .I(dataWriteZ0Z_4));
    InMux I__8546 (
            .O(N__36384),
            .I(N__36381));
    LocalMux I__8545 (
            .O(N__36381),
            .I(\PWMInstance2.PWMPulseWidthCountZ0Z_4 ));
    CascadeMux I__8544 (
            .O(N__36378),
            .I(N__36373));
    InMux I__8543 (
            .O(N__36377),
            .I(N__36363));
    InMux I__8542 (
            .O(N__36376),
            .I(N__36359));
    InMux I__8541 (
            .O(N__36373),
            .I(N__36348));
    InMux I__8540 (
            .O(N__36372),
            .I(N__36348));
    InMux I__8539 (
            .O(N__36371),
            .I(N__36348));
    InMux I__8538 (
            .O(N__36370),
            .I(N__36348));
    InMux I__8537 (
            .O(N__36369),
            .I(N__36348));
    InMux I__8536 (
            .O(N__36368),
            .I(N__36342));
    InMux I__8535 (
            .O(N__36367),
            .I(N__36339));
    InMux I__8534 (
            .O(N__36366),
            .I(N__36336));
    LocalMux I__8533 (
            .O(N__36363),
            .I(N__36333));
    InMux I__8532 (
            .O(N__36362),
            .I(N__36329));
    LocalMux I__8531 (
            .O(N__36359),
            .I(N__36326));
    LocalMux I__8530 (
            .O(N__36348),
            .I(N__36323));
    InMux I__8529 (
            .O(N__36347),
            .I(N__36320));
    InMux I__8528 (
            .O(N__36346),
            .I(N__36317));
    InMux I__8527 (
            .O(N__36345),
            .I(N__36314));
    LocalMux I__8526 (
            .O(N__36342),
            .I(N__36311));
    LocalMux I__8525 (
            .O(N__36339),
            .I(N__36308));
    LocalMux I__8524 (
            .O(N__36336),
            .I(N__36305));
    Span4Mux_v I__8523 (
            .O(N__36333),
            .I(N__36302));
    InMux I__8522 (
            .O(N__36332),
            .I(N__36299));
    LocalMux I__8521 (
            .O(N__36329),
            .I(N__36296));
    Span4Mux_v I__8520 (
            .O(N__36326),
            .I(N__36293));
    Span4Mux_v I__8519 (
            .O(N__36323),
            .I(N__36290));
    LocalMux I__8518 (
            .O(N__36320),
            .I(N__36285));
    LocalMux I__8517 (
            .O(N__36317),
            .I(N__36285));
    LocalMux I__8516 (
            .O(N__36314),
            .I(N__36281));
    Span4Mux_v I__8515 (
            .O(N__36311),
            .I(N__36278));
    Span4Mux_v I__8514 (
            .O(N__36308),
            .I(N__36271));
    Span4Mux_v I__8513 (
            .O(N__36305),
            .I(N__36271));
    Span4Mux_v I__8512 (
            .O(N__36302),
            .I(N__36271));
    LocalMux I__8511 (
            .O(N__36299),
            .I(N__36266));
    Span4Mux_v I__8510 (
            .O(N__36296),
            .I(N__36266));
    Span4Mux_h I__8509 (
            .O(N__36293),
            .I(N__36263));
    Span4Mux_h I__8508 (
            .O(N__36290),
            .I(N__36260));
    Span4Mux_h I__8507 (
            .O(N__36285),
            .I(N__36257));
    InMux I__8506 (
            .O(N__36284),
            .I(N__36254));
    Span4Mux_h I__8505 (
            .O(N__36281),
            .I(N__36251));
    Span4Mux_v I__8504 (
            .O(N__36278),
            .I(N__36246));
    Span4Mux_h I__8503 (
            .O(N__36271),
            .I(N__36246));
    Span4Mux_v I__8502 (
            .O(N__36266),
            .I(N__36239));
    Span4Mux_h I__8501 (
            .O(N__36263),
            .I(N__36239));
    Span4Mux_v I__8500 (
            .O(N__36260),
            .I(N__36239));
    Span4Mux_v I__8499 (
            .O(N__36257),
            .I(N__36236));
    LocalMux I__8498 (
            .O(N__36254),
            .I(dataWriteZ0Z_5));
    Odrv4 I__8497 (
            .O(N__36251),
            .I(dataWriteZ0Z_5));
    Odrv4 I__8496 (
            .O(N__36246),
            .I(dataWriteZ0Z_5));
    Odrv4 I__8495 (
            .O(N__36239),
            .I(dataWriteZ0Z_5));
    Odrv4 I__8494 (
            .O(N__36236),
            .I(dataWriteZ0Z_5));
    InMux I__8493 (
            .O(N__36225),
            .I(N__36222));
    LocalMux I__8492 (
            .O(N__36222),
            .I(\PWMInstance2.PWMPulseWidthCountZ0Z_5 ));
    InMux I__8491 (
            .O(N__36219),
            .I(N__36212));
    InMux I__8490 (
            .O(N__36218),
            .I(N__36212));
    InMux I__8489 (
            .O(N__36217),
            .I(N__36209));
    LocalMux I__8488 (
            .O(N__36212),
            .I(N__36206));
    LocalMux I__8487 (
            .O(N__36209),
            .I(\PWMInstance2.periodCounterZ0Z_10 ));
    Odrv4 I__8486 (
            .O(N__36206),
            .I(\PWMInstance2.periodCounterZ0Z_10 ));
    CascadeMux I__8485 (
            .O(N__36201),
            .I(N__36197));
    CascadeMux I__8484 (
            .O(N__36200),
            .I(N__36193));
    InMux I__8483 (
            .O(N__36197),
            .I(N__36190));
    InMux I__8482 (
            .O(N__36196),
            .I(N__36187));
    InMux I__8481 (
            .O(N__36193),
            .I(N__36184));
    LocalMux I__8480 (
            .O(N__36190),
            .I(N__36181));
    LocalMux I__8479 (
            .O(N__36187),
            .I(\PWMInstance2.periodCounterZ0Z_11 ));
    LocalMux I__8478 (
            .O(N__36184),
            .I(\PWMInstance2.periodCounterZ0Z_11 ));
    Odrv4 I__8477 (
            .O(N__36181),
            .I(\PWMInstance2.periodCounterZ0Z_11 ));
    InMux I__8476 (
            .O(N__36174),
            .I(N__36171));
    LocalMux I__8475 (
            .O(N__36171),
            .I(\PWMInstance2.un1_PWMPulseWidthCount_0_I_33_c_RNO_1 ));
    InMux I__8474 (
            .O(N__36168),
            .I(N__36161));
    InMux I__8473 (
            .O(N__36167),
            .I(N__36154));
    InMux I__8472 (
            .O(N__36166),
            .I(N__36151));
    InMux I__8471 (
            .O(N__36165),
            .I(N__36146));
    CascadeMux I__8470 (
            .O(N__36164),
            .I(N__36143));
    LocalMux I__8469 (
            .O(N__36161),
            .I(N__36139));
    InMux I__8468 (
            .O(N__36160),
            .I(N__36136));
    InMux I__8467 (
            .O(N__36159),
            .I(N__36130));
    InMux I__8466 (
            .O(N__36158),
            .I(N__36127));
    InMux I__8465 (
            .O(N__36157),
            .I(N__36124));
    LocalMux I__8464 (
            .O(N__36154),
            .I(N__36121));
    LocalMux I__8463 (
            .O(N__36151),
            .I(N__36118));
    InMux I__8462 (
            .O(N__36150),
            .I(N__36115));
    InMux I__8461 (
            .O(N__36149),
            .I(N__36112));
    LocalMux I__8460 (
            .O(N__36146),
            .I(N__36109));
    InMux I__8459 (
            .O(N__36143),
            .I(N__36106));
    InMux I__8458 (
            .O(N__36142),
            .I(N__36103));
    Span4Mux_v I__8457 (
            .O(N__36139),
            .I(N__36098));
    LocalMux I__8456 (
            .O(N__36136),
            .I(N__36098));
    InMux I__8455 (
            .O(N__36135),
            .I(N__36095));
    InMux I__8454 (
            .O(N__36134),
            .I(N__36090));
    InMux I__8453 (
            .O(N__36133),
            .I(N__36090));
    LocalMux I__8452 (
            .O(N__36130),
            .I(N__36084));
    LocalMux I__8451 (
            .O(N__36127),
            .I(N__36084));
    LocalMux I__8450 (
            .O(N__36124),
            .I(N__36081));
    Span4Mux_v I__8449 (
            .O(N__36121),
            .I(N__36076));
    Span4Mux_v I__8448 (
            .O(N__36118),
            .I(N__36076));
    LocalMux I__8447 (
            .O(N__36115),
            .I(N__36073));
    LocalMux I__8446 (
            .O(N__36112),
            .I(N__36070));
    Sp12to4 I__8445 (
            .O(N__36109),
            .I(N__36065));
    LocalMux I__8444 (
            .O(N__36106),
            .I(N__36065));
    LocalMux I__8443 (
            .O(N__36103),
            .I(N__36062));
    Span4Mux_h I__8442 (
            .O(N__36098),
            .I(N__36055));
    LocalMux I__8441 (
            .O(N__36095),
            .I(N__36055));
    LocalMux I__8440 (
            .O(N__36090),
            .I(N__36055));
    InMux I__8439 (
            .O(N__36089),
            .I(N__36052));
    Span4Mux_v I__8438 (
            .O(N__36084),
            .I(N__36049));
    Span4Mux_h I__8437 (
            .O(N__36081),
            .I(N__36046));
    Sp12to4 I__8436 (
            .O(N__36076),
            .I(N__36037));
    Span12Mux_s9_v I__8435 (
            .O(N__36073),
            .I(N__36037));
    Span12Mux_s6_h I__8434 (
            .O(N__36070),
            .I(N__36037));
    Span12Mux_s10_v I__8433 (
            .O(N__36065),
            .I(N__36037));
    Span4Mux_h I__8432 (
            .O(N__36062),
            .I(N__36030));
    Span4Mux_h I__8431 (
            .O(N__36055),
            .I(N__36030));
    LocalMux I__8430 (
            .O(N__36052),
            .I(N__36030));
    Odrv4 I__8429 (
            .O(N__36049),
            .I(dataWriteZ0Z_10));
    Odrv4 I__8428 (
            .O(N__36046),
            .I(dataWriteZ0Z_10));
    Odrv12 I__8427 (
            .O(N__36037),
            .I(dataWriteZ0Z_10));
    Odrv4 I__8426 (
            .O(N__36030),
            .I(dataWriteZ0Z_10));
    InMux I__8425 (
            .O(N__36021),
            .I(N__36018));
    LocalMux I__8424 (
            .O(N__36018),
            .I(\PWMInstance2.PWMPulseWidthCountZ0Z_10 ));
    CascadeMux I__8423 (
            .O(N__36015),
            .I(N__36007));
    InMux I__8422 (
            .O(N__36014),
            .I(N__35999));
    InMux I__8421 (
            .O(N__36013),
            .I(N__35995));
    InMux I__8420 (
            .O(N__36012),
            .I(N__35990));
    InMux I__8419 (
            .O(N__36011),
            .I(N__35987));
    InMux I__8418 (
            .O(N__36010),
            .I(N__35978));
    InMux I__8417 (
            .O(N__36007),
            .I(N__35978));
    InMux I__8416 (
            .O(N__36006),
            .I(N__35978));
    InMux I__8415 (
            .O(N__36005),
            .I(N__35978));
    InMux I__8414 (
            .O(N__36004),
            .I(N__35975));
    InMux I__8413 (
            .O(N__36003),
            .I(N__35970));
    InMux I__8412 (
            .O(N__36002),
            .I(N__35967));
    LocalMux I__8411 (
            .O(N__35999),
            .I(N__35964));
    InMux I__8410 (
            .O(N__35998),
            .I(N__35961));
    LocalMux I__8409 (
            .O(N__35995),
            .I(N__35958));
    InMux I__8408 (
            .O(N__35994),
            .I(N__35955));
    InMux I__8407 (
            .O(N__35993),
            .I(N__35952));
    LocalMux I__8406 (
            .O(N__35990),
            .I(N__35949));
    LocalMux I__8405 (
            .O(N__35987),
            .I(N__35944));
    LocalMux I__8404 (
            .O(N__35978),
            .I(N__35944));
    LocalMux I__8403 (
            .O(N__35975),
            .I(N__35941));
    InMux I__8402 (
            .O(N__35974),
            .I(N__35938));
    CascadeMux I__8401 (
            .O(N__35973),
            .I(N__35935));
    LocalMux I__8400 (
            .O(N__35970),
            .I(N__35930));
    LocalMux I__8399 (
            .O(N__35967),
            .I(N__35930));
    Span4Mux_v I__8398 (
            .O(N__35964),
            .I(N__35927));
    LocalMux I__8397 (
            .O(N__35961),
            .I(N__35924));
    Span4Mux_h I__8396 (
            .O(N__35958),
            .I(N__35919));
    LocalMux I__8395 (
            .O(N__35955),
            .I(N__35919));
    LocalMux I__8394 (
            .O(N__35952),
            .I(N__35916));
    Span4Mux_v I__8393 (
            .O(N__35949),
            .I(N__35911));
    Span4Mux_h I__8392 (
            .O(N__35944),
            .I(N__35911));
    Span4Mux_h I__8391 (
            .O(N__35941),
            .I(N__35906));
    LocalMux I__8390 (
            .O(N__35938),
            .I(N__35906));
    InMux I__8389 (
            .O(N__35935),
            .I(N__35903));
    Span12Mux_s10_v I__8388 (
            .O(N__35930),
            .I(N__35900));
    Span4Mux_v I__8387 (
            .O(N__35927),
            .I(N__35897));
    Span4Mux_h I__8386 (
            .O(N__35924),
            .I(N__35892));
    Span4Mux_h I__8385 (
            .O(N__35919),
            .I(N__35892));
    Span4Mux_v I__8384 (
            .O(N__35916),
            .I(N__35887));
    Span4Mux_h I__8383 (
            .O(N__35911),
            .I(N__35887));
    Span4Mux_h I__8382 (
            .O(N__35906),
            .I(N__35882));
    LocalMux I__8381 (
            .O(N__35903),
            .I(N__35882));
    Odrv12 I__8380 (
            .O(N__35900),
            .I(dataWriteZ0Z_11));
    Odrv4 I__8379 (
            .O(N__35897),
            .I(dataWriteZ0Z_11));
    Odrv4 I__8378 (
            .O(N__35892),
            .I(dataWriteZ0Z_11));
    Odrv4 I__8377 (
            .O(N__35887),
            .I(dataWriteZ0Z_11));
    Odrv4 I__8376 (
            .O(N__35882),
            .I(dataWriteZ0Z_11));
    InMux I__8375 (
            .O(N__35871),
            .I(N__35868));
    LocalMux I__8374 (
            .O(N__35868),
            .I(\PWMInstance2.PWMPulseWidthCountZ0Z_11 ));
    CEMux I__8373 (
            .O(N__35865),
            .I(N__35862));
    LocalMux I__8372 (
            .O(N__35862),
            .I(N__35858));
    CEMux I__8371 (
            .O(N__35861),
            .I(N__35855));
    Span4Mux_v I__8370 (
            .O(N__35858),
            .I(N__35848));
    LocalMux I__8369 (
            .O(N__35855),
            .I(N__35848));
    CEMux I__8368 (
            .O(N__35854),
            .I(N__35845));
    CEMux I__8367 (
            .O(N__35853),
            .I(N__35842));
    Span4Mux_h I__8366 (
            .O(N__35848),
            .I(N__35839));
    LocalMux I__8365 (
            .O(N__35845),
            .I(\PWMInstance2.pwmWrite_0_2 ));
    LocalMux I__8364 (
            .O(N__35842),
            .I(\PWMInstance2.pwmWrite_0_2 ));
    Odrv4 I__8363 (
            .O(N__35839),
            .I(\PWMInstance2.pwmWrite_0_2 ));
    InMux I__8362 (
            .O(N__35832),
            .I(N__35821));
    InMux I__8361 (
            .O(N__35831),
            .I(N__35818));
    InMux I__8360 (
            .O(N__35830),
            .I(N__35815));
    InMux I__8359 (
            .O(N__35829),
            .I(N__35812));
    InMux I__8358 (
            .O(N__35828),
            .I(N__35809));
    InMux I__8357 (
            .O(N__35827),
            .I(N__35806));
    InMux I__8356 (
            .O(N__35826),
            .I(N__35803));
    InMux I__8355 (
            .O(N__35825),
            .I(N__35800));
    InMux I__8354 (
            .O(N__35824),
            .I(N__35797));
    LocalMux I__8353 (
            .O(N__35821),
            .I(N__35790));
    LocalMux I__8352 (
            .O(N__35818),
            .I(N__35778));
    LocalMux I__8351 (
            .O(N__35815),
            .I(N__35766));
    LocalMux I__8350 (
            .O(N__35812),
            .I(N__35760));
    LocalMux I__8349 (
            .O(N__35809),
            .I(N__35749));
    LocalMux I__8348 (
            .O(N__35806),
            .I(N__35744));
    LocalMux I__8347 (
            .O(N__35803),
            .I(N__35730));
    LocalMux I__8346 (
            .O(N__35800),
            .I(N__35710));
    LocalMux I__8345 (
            .O(N__35797),
            .I(N__35686));
    SRMux I__8344 (
            .O(N__35796),
            .I(N__35469));
    SRMux I__8343 (
            .O(N__35795),
            .I(N__35469));
    SRMux I__8342 (
            .O(N__35794),
            .I(N__35469));
    SRMux I__8341 (
            .O(N__35793),
            .I(N__35469));
    Glb2LocalMux I__8340 (
            .O(N__35790),
            .I(N__35469));
    SRMux I__8339 (
            .O(N__35789),
            .I(N__35469));
    SRMux I__8338 (
            .O(N__35788),
            .I(N__35469));
    SRMux I__8337 (
            .O(N__35787),
            .I(N__35469));
    SRMux I__8336 (
            .O(N__35786),
            .I(N__35469));
    SRMux I__8335 (
            .O(N__35785),
            .I(N__35469));
    SRMux I__8334 (
            .O(N__35784),
            .I(N__35469));
    SRMux I__8333 (
            .O(N__35783),
            .I(N__35469));
    SRMux I__8332 (
            .O(N__35782),
            .I(N__35469));
    SRMux I__8331 (
            .O(N__35781),
            .I(N__35469));
    Glb2LocalMux I__8330 (
            .O(N__35778),
            .I(N__35469));
    SRMux I__8329 (
            .O(N__35777),
            .I(N__35469));
    SRMux I__8328 (
            .O(N__35776),
            .I(N__35469));
    SRMux I__8327 (
            .O(N__35775),
            .I(N__35469));
    SRMux I__8326 (
            .O(N__35774),
            .I(N__35469));
    SRMux I__8325 (
            .O(N__35773),
            .I(N__35469));
    SRMux I__8324 (
            .O(N__35772),
            .I(N__35469));
    SRMux I__8323 (
            .O(N__35771),
            .I(N__35469));
    SRMux I__8322 (
            .O(N__35770),
            .I(N__35469));
    SRMux I__8321 (
            .O(N__35769),
            .I(N__35469));
    Glb2LocalMux I__8320 (
            .O(N__35766),
            .I(N__35469));
    SRMux I__8319 (
            .O(N__35765),
            .I(N__35469));
    SRMux I__8318 (
            .O(N__35764),
            .I(N__35469));
    SRMux I__8317 (
            .O(N__35763),
            .I(N__35469));
    Glb2LocalMux I__8316 (
            .O(N__35760),
            .I(N__35469));
    SRMux I__8315 (
            .O(N__35759),
            .I(N__35469));
    SRMux I__8314 (
            .O(N__35758),
            .I(N__35469));
    SRMux I__8313 (
            .O(N__35757),
            .I(N__35469));
    SRMux I__8312 (
            .O(N__35756),
            .I(N__35469));
    SRMux I__8311 (
            .O(N__35755),
            .I(N__35469));
    SRMux I__8310 (
            .O(N__35754),
            .I(N__35469));
    SRMux I__8309 (
            .O(N__35753),
            .I(N__35469));
    SRMux I__8308 (
            .O(N__35752),
            .I(N__35469));
    Glb2LocalMux I__8307 (
            .O(N__35749),
            .I(N__35469));
    SRMux I__8306 (
            .O(N__35748),
            .I(N__35469));
    SRMux I__8305 (
            .O(N__35747),
            .I(N__35469));
    Glb2LocalMux I__8304 (
            .O(N__35744),
            .I(N__35469));
    SRMux I__8303 (
            .O(N__35743),
            .I(N__35469));
    SRMux I__8302 (
            .O(N__35742),
            .I(N__35469));
    SRMux I__8301 (
            .O(N__35741),
            .I(N__35469));
    SRMux I__8300 (
            .O(N__35740),
            .I(N__35469));
    SRMux I__8299 (
            .O(N__35739),
            .I(N__35469));
    SRMux I__8298 (
            .O(N__35738),
            .I(N__35469));
    SRMux I__8297 (
            .O(N__35737),
            .I(N__35469));
    SRMux I__8296 (
            .O(N__35736),
            .I(N__35469));
    SRMux I__8295 (
            .O(N__35735),
            .I(N__35469));
    SRMux I__8294 (
            .O(N__35734),
            .I(N__35469));
    SRMux I__8293 (
            .O(N__35733),
            .I(N__35469));
    Glb2LocalMux I__8292 (
            .O(N__35730),
            .I(N__35469));
    SRMux I__8291 (
            .O(N__35729),
            .I(N__35469));
    SRMux I__8290 (
            .O(N__35728),
            .I(N__35469));
    SRMux I__8289 (
            .O(N__35727),
            .I(N__35469));
    SRMux I__8288 (
            .O(N__35726),
            .I(N__35469));
    SRMux I__8287 (
            .O(N__35725),
            .I(N__35469));
    SRMux I__8286 (
            .O(N__35724),
            .I(N__35469));
    SRMux I__8285 (
            .O(N__35723),
            .I(N__35469));
    SRMux I__8284 (
            .O(N__35722),
            .I(N__35469));
    SRMux I__8283 (
            .O(N__35721),
            .I(N__35469));
    SRMux I__8282 (
            .O(N__35720),
            .I(N__35469));
    SRMux I__8281 (
            .O(N__35719),
            .I(N__35469));
    SRMux I__8280 (
            .O(N__35718),
            .I(N__35469));
    SRMux I__8279 (
            .O(N__35717),
            .I(N__35469));
    SRMux I__8278 (
            .O(N__35716),
            .I(N__35469));
    SRMux I__8277 (
            .O(N__35715),
            .I(N__35469));
    SRMux I__8276 (
            .O(N__35714),
            .I(N__35469));
    SRMux I__8275 (
            .O(N__35713),
            .I(N__35469));
    Glb2LocalMux I__8274 (
            .O(N__35710),
            .I(N__35469));
    SRMux I__8273 (
            .O(N__35709),
            .I(N__35469));
    SRMux I__8272 (
            .O(N__35708),
            .I(N__35469));
    SRMux I__8271 (
            .O(N__35707),
            .I(N__35469));
    SRMux I__8270 (
            .O(N__35706),
            .I(N__35469));
    SRMux I__8269 (
            .O(N__35705),
            .I(N__35469));
    SRMux I__8268 (
            .O(N__35704),
            .I(N__35469));
    SRMux I__8267 (
            .O(N__35703),
            .I(N__35469));
    SRMux I__8266 (
            .O(N__35702),
            .I(N__35469));
    SRMux I__8265 (
            .O(N__35701),
            .I(N__35469));
    SRMux I__8264 (
            .O(N__35700),
            .I(N__35469));
    SRMux I__8263 (
            .O(N__35699),
            .I(N__35469));
    SRMux I__8262 (
            .O(N__35698),
            .I(N__35469));
    SRMux I__8261 (
            .O(N__35697),
            .I(N__35469));
    SRMux I__8260 (
            .O(N__35696),
            .I(N__35469));
    SRMux I__8259 (
            .O(N__35695),
            .I(N__35469));
    SRMux I__8258 (
            .O(N__35694),
            .I(N__35469));
    SRMux I__8257 (
            .O(N__35693),
            .I(N__35469));
    SRMux I__8256 (
            .O(N__35692),
            .I(N__35469));
    SRMux I__8255 (
            .O(N__35691),
            .I(N__35469));
    SRMux I__8254 (
            .O(N__35690),
            .I(N__35469));
    SRMux I__8253 (
            .O(N__35689),
            .I(N__35469));
    Glb2LocalMux I__8252 (
            .O(N__35686),
            .I(N__35469));
    SRMux I__8251 (
            .O(N__35685),
            .I(N__35469));
    SRMux I__8250 (
            .O(N__35684),
            .I(N__35469));
    SRMux I__8249 (
            .O(N__35683),
            .I(N__35469));
    SRMux I__8248 (
            .O(N__35682),
            .I(N__35469));
    SRMux I__8247 (
            .O(N__35681),
            .I(N__35469));
    SRMux I__8246 (
            .O(N__35680),
            .I(N__35469));
    SRMux I__8245 (
            .O(N__35679),
            .I(N__35469));
    SRMux I__8244 (
            .O(N__35678),
            .I(N__35469));
    SRMux I__8243 (
            .O(N__35677),
            .I(N__35469));
    SRMux I__8242 (
            .O(N__35676),
            .I(N__35469));
    GlobalMux I__8241 (
            .O(N__35469),
            .I(N__35466));
    gio2CtrlBuf I__8240 (
            .O(N__35466),
            .I(RST_c_i_g));
    IoInMux I__8239 (
            .O(N__35463),
            .I(N__35460));
    LocalMux I__8238 (
            .O(N__35460),
            .I(PWM2_obufLegalizeSB_DFFNet));
    InMux I__8237 (
            .O(N__35457),
            .I(N__35452));
    InMux I__8236 (
            .O(N__35456),
            .I(N__35449));
    InMux I__8235 (
            .O(N__35455),
            .I(N__35446));
    LocalMux I__8234 (
            .O(N__35452),
            .I(\PWMInstance2.periodCounterZ0Z_9 ));
    LocalMux I__8233 (
            .O(N__35449),
            .I(\PWMInstance2.periodCounterZ0Z_9 ));
    LocalMux I__8232 (
            .O(N__35446),
            .I(\PWMInstance2.periodCounterZ0Z_9 ));
    InMux I__8231 (
            .O(N__35439),
            .I(\PWMInstance2.un1_periodCounter_2_cry_8 ));
    InMux I__8230 (
            .O(N__35436),
            .I(\PWMInstance2.un1_periodCounter_2_cry_9 ));
    InMux I__8229 (
            .O(N__35433),
            .I(\PWMInstance2.un1_periodCounter_2_cry_10 ));
    InMux I__8228 (
            .O(N__35430),
            .I(\PWMInstance2.un1_periodCounter_2_cry_11 ));
    CascadeMux I__8227 (
            .O(N__35427),
            .I(N__35423));
    InMux I__8226 (
            .O(N__35426),
            .I(N__35419));
    InMux I__8225 (
            .O(N__35423),
            .I(N__35416));
    InMux I__8224 (
            .O(N__35422),
            .I(N__35413));
    LocalMux I__8223 (
            .O(N__35419),
            .I(\PWMInstance2.periodCounterZ0Z_13 ));
    LocalMux I__8222 (
            .O(N__35416),
            .I(\PWMInstance2.periodCounterZ0Z_13 ));
    LocalMux I__8221 (
            .O(N__35413),
            .I(\PWMInstance2.periodCounterZ0Z_13 ));
    InMux I__8220 (
            .O(N__35406),
            .I(\PWMInstance2.un1_periodCounter_2_cry_12 ));
    InMux I__8219 (
            .O(N__35403),
            .I(\PWMInstance2.un1_periodCounter_2_cry_13 ));
    CascadeMux I__8218 (
            .O(N__35400),
            .I(N__35396));
    InMux I__8217 (
            .O(N__35399),
            .I(N__35392));
    InMux I__8216 (
            .O(N__35396),
            .I(N__35389));
    InMux I__8215 (
            .O(N__35395),
            .I(N__35386));
    LocalMux I__8214 (
            .O(N__35392),
            .I(\PWMInstance2.periodCounterZ0Z_15 ));
    LocalMux I__8213 (
            .O(N__35389),
            .I(\PWMInstance2.periodCounterZ0Z_15 ));
    LocalMux I__8212 (
            .O(N__35386),
            .I(\PWMInstance2.periodCounterZ0Z_15 ));
    InMux I__8211 (
            .O(N__35379),
            .I(\PWMInstance2.un1_periodCounter_2_cry_14 ));
    CascadeMux I__8210 (
            .O(N__35376),
            .I(N__35373));
    InMux I__8209 (
            .O(N__35373),
            .I(N__35365));
    InMux I__8208 (
            .O(N__35372),
            .I(N__35362));
    InMux I__8207 (
            .O(N__35371),
            .I(N__35359));
    InMux I__8206 (
            .O(N__35370),
            .I(N__35354));
    InMux I__8205 (
            .O(N__35369),
            .I(N__35354));
    InMux I__8204 (
            .O(N__35368),
            .I(N__35351));
    LocalMux I__8203 (
            .O(N__35365),
            .I(N__35348));
    LocalMux I__8202 (
            .O(N__35362),
            .I(\PWMInstance2.out_0_sqmuxa ));
    LocalMux I__8201 (
            .O(N__35359),
            .I(\PWMInstance2.out_0_sqmuxa ));
    LocalMux I__8200 (
            .O(N__35354),
            .I(\PWMInstance2.out_0_sqmuxa ));
    LocalMux I__8199 (
            .O(N__35351),
            .I(\PWMInstance2.out_0_sqmuxa ));
    Odrv4 I__8198 (
            .O(N__35348),
            .I(\PWMInstance2.out_0_sqmuxa ));
    InMux I__8197 (
            .O(N__35337),
            .I(bfn_18_13_0_));
    CascadeMux I__8196 (
            .O(N__35334),
            .I(N__35330));
    InMux I__8195 (
            .O(N__35333),
            .I(N__35326));
    InMux I__8194 (
            .O(N__35330),
            .I(N__35321));
    InMux I__8193 (
            .O(N__35329),
            .I(N__35321));
    LocalMux I__8192 (
            .O(N__35326),
            .I(\PWMInstance2.periodCounterZ0Z_16 ));
    LocalMux I__8191 (
            .O(N__35321),
            .I(\PWMInstance2.periodCounterZ0Z_16 ));
    SRMux I__8190 (
            .O(N__35316),
            .I(N__35244));
    SRMux I__8189 (
            .O(N__35315),
            .I(N__35244));
    SRMux I__8188 (
            .O(N__35314),
            .I(N__35244));
    SRMux I__8187 (
            .O(N__35313),
            .I(N__35244));
    SRMux I__8186 (
            .O(N__35312),
            .I(N__35244));
    SRMux I__8185 (
            .O(N__35311),
            .I(N__35244));
    SRMux I__8184 (
            .O(N__35310),
            .I(N__35244));
    SRMux I__8183 (
            .O(N__35309),
            .I(N__35244));
    SRMux I__8182 (
            .O(N__35308),
            .I(N__35244));
    SRMux I__8181 (
            .O(N__35307),
            .I(N__35244));
    SRMux I__8180 (
            .O(N__35306),
            .I(N__35244));
    SRMux I__8179 (
            .O(N__35305),
            .I(N__35244));
    SRMux I__8178 (
            .O(N__35304),
            .I(N__35244));
    SRMux I__8177 (
            .O(N__35303),
            .I(N__35244));
    SRMux I__8176 (
            .O(N__35302),
            .I(N__35244));
    SRMux I__8175 (
            .O(N__35301),
            .I(N__35244));
    SRMux I__8174 (
            .O(N__35300),
            .I(N__35244));
    SRMux I__8173 (
            .O(N__35299),
            .I(N__35244));
    SRMux I__8172 (
            .O(N__35298),
            .I(N__35244));
    SRMux I__8171 (
            .O(N__35297),
            .I(N__35244));
    SRMux I__8170 (
            .O(N__35296),
            .I(N__35244));
    SRMux I__8169 (
            .O(N__35295),
            .I(N__35244));
    SRMux I__8168 (
            .O(N__35294),
            .I(N__35244));
    SRMux I__8167 (
            .O(N__35293),
            .I(N__35244));
    GlobalMux I__8166 (
            .O(N__35244),
            .I(N__35241));
    gio2CtrlBuf I__8165 (
            .O(N__35241),
            .I(PWMInstance0_N_42_g));
    CascadeMux I__8164 (
            .O(N__35238),
            .I(N__35234));
    InMux I__8163 (
            .O(N__35237),
            .I(N__35230));
    InMux I__8162 (
            .O(N__35234),
            .I(N__35227));
    InMux I__8161 (
            .O(N__35233),
            .I(N__35224));
    LocalMux I__8160 (
            .O(N__35230),
            .I(N__35219));
    LocalMux I__8159 (
            .O(N__35227),
            .I(N__35219));
    LocalMux I__8158 (
            .O(N__35224),
            .I(\PWMInstance2.periodCounterZ0Z_5 ));
    Odrv4 I__8157 (
            .O(N__35219),
            .I(\PWMInstance2.periodCounterZ0Z_5 ));
    InMux I__8156 (
            .O(N__35214),
            .I(N__35211));
    LocalMux I__8155 (
            .O(N__35211),
            .I(\PWMInstance2.un1_PWMPulseWidthCount_0_I_15_c_RNO_1 ));
    CascadeMux I__8154 (
            .O(N__35208),
            .I(N__35203));
    InMux I__8153 (
            .O(N__35207),
            .I(N__35200));
    InMux I__8152 (
            .O(N__35206),
            .I(N__35197));
    InMux I__8151 (
            .O(N__35203),
            .I(N__35194));
    LocalMux I__8150 (
            .O(N__35200),
            .I(\PWMInstance2.periodCounterZ0Z_1 ));
    LocalMux I__8149 (
            .O(N__35197),
            .I(\PWMInstance2.periodCounterZ0Z_1 ));
    LocalMux I__8148 (
            .O(N__35194),
            .I(\PWMInstance2.periodCounterZ0Z_1 ));
    InMux I__8147 (
            .O(N__35187),
            .I(\PWMInstance2.un1_periodCounter_2_cry_0 ));
    InMux I__8146 (
            .O(N__35184),
            .I(\PWMInstance2.un1_periodCounter_2_cry_1 ));
    InMux I__8145 (
            .O(N__35181),
            .I(N__35174));
    InMux I__8144 (
            .O(N__35180),
            .I(N__35174));
    InMux I__8143 (
            .O(N__35179),
            .I(N__35171));
    LocalMux I__8142 (
            .O(N__35174),
            .I(N__35168));
    LocalMux I__8141 (
            .O(N__35171),
            .I(\PWMInstance2.periodCounterZ0Z_3 ));
    Odrv4 I__8140 (
            .O(N__35168),
            .I(\PWMInstance2.periodCounterZ0Z_3 ));
    InMux I__8139 (
            .O(N__35163),
            .I(\PWMInstance2.un1_periodCounter_2_cry_2 ));
    InMux I__8138 (
            .O(N__35160),
            .I(\PWMInstance2.un1_periodCounter_2_cry_3 ));
    InMux I__8137 (
            .O(N__35157),
            .I(\PWMInstance2.un1_periodCounter_2_cry_4 ));
    CascadeMux I__8136 (
            .O(N__35154),
            .I(N__35149));
    CascadeMux I__8135 (
            .O(N__35153),
            .I(N__35146));
    InMux I__8134 (
            .O(N__35152),
            .I(N__35143));
    InMux I__8133 (
            .O(N__35149),
            .I(N__35138));
    InMux I__8132 (
            .O(N__35146),
            .I(N__35138));
    LocalMux I__8131 (
            .O(N__35143),
            .I(\PWMInstance2.periodCounterZ0Z_6 ));
    LocalMux I__8130 (
            .O(N__35138),
            .I(\PWMInstance2.periodCounterZ0Z_6 ));
    InMux I__8129 (
            .O(N__35133),
            .I(\PWMInstance2.un1_periodCounter_2_cry_5 ));
    InMux I__8128 (
            .O(N__35130),
            .I(N__35125));
    InMux I__8127 (
            .O(N__35129),
            .I(N__35122));
    InMux I__8126 (
            .O(N__35128),
            .I(N__35119));
    LocalMux I__8125 (
            .O(N__35125),
            .I(\PWMInstance2.periodCounterZ0Z_7 ));
    LocalMux I__8124 (
            .O(N__35122),
            .I(\PWMInstance2.periodCounterZ0Z_7 ));
    LocalMux I__8123 (
            .O(N__35119),
            .I(\PWMInstance2.periodCounterZ0Z_7 ));
    InMux I__8122 (
            .O(N__35112),
            .I(\PWMInstance2.un1_periodCounter_2_cry_6 ));
    CascadeMux I__8121 (
            .O(N__35109),
            .I(N__35104));
    InMux I__8120 (
            .O(N__35108),
            .I(N__35101));
    InMux I__8119 (
            .O(N__35107),
            .I(N__35096));
    InMux I__8118 (
            .O(N__35104),
            .I(N__35096));
    LocalMux I__8117 (
            .O(N__35101),
            .I(\PWMInstance2.periodCounterZ0Z_8 ));
    LocalMux I__8116 (
            .O(N__35096),
            .I(\PWMInstance2.periodCounterZ0Z_8 ));
    InMux I__8115 (
            .O(N__35091),
            .I(bfn_18_12_0_));
    InMux I__8114 (
            .O(N__35088),
            .I(N__35076));
    InMux I__8113 (
            .O(N__35087),
            .I(N__35076));
    InMux I__8112 (
            .O(N__35086),
            .I(N__35076));
    InMux I__8111 (
            .O(N__35085),
            .I(N__35076));
    LocalMux I__8110 (
            .O(N__35076),
            .I(N__35073));
    Span4Mux_v I__8109 (
            .O(N__35073),
            .I(N__35070));
    Span4Mux_h I__8108 (
            .O(N__35070),
            .I(N__35067));
    Span4Mux_h I__8107 (
            .O(N__35067),
            .I(N__35064));
    Odrv4 I__8106 (
            .O(N__35064),
            .I(MOSIrZ0Z_1));
    InMux I__8105 (
            .O(N__35061),
            .I(N__35057));
    InMux I__8104 (
            .O(N__35060),
            .I(N__35054));
    LocalMux I__8103 (
            .O(N__35057),
            .I(N__35051));
    LocalMux I__8102 (
            .O(N__35054),
            .I(N__35047));
    Span4Mux_v I__8101 (
            .O(N__35051),
            .I(N__35044));
    InMux I__8100 (
            .O(N__35050),
            .I(N__35041));
    Span4Mux_h I__8099 (
            .O(N__35047),
            .I(N__35038));
    Span4Mux_v I__8098 (
            .O(N__35044),
            .I(N__35033));
    LocalMux I__8097 (
            .O(N__35041),
            .I(N__35033));
    Span4Mux_h I__8096 (
            .O(N__35038),
            .I(N__35030));
    Odrv4 I__8095 (
            .O(N__35033),
            .I(dataRead1_10));
    Odrv4 I__8094 (
            .O(N__35030),
            .I(dataRead1_10));
    CascadeMux I__8093 (
            .O(N__35025),
            .I(N__35021));
    CascadeMux I__8092 (
            .O(N__35024),
            .I(N__35018));
    InMux I__8091 (
            .O(N__35021),
            .I(N__35015));
    InMux I__8090 (
            .O(N__35018),
            .I(N__35012));
    LocalMux I__8089 (
            .O(N__35015),
            .I(N__35009));
    LocalMux I__8088 (
            .O(N__35012),
            .I(N__35005));
    Span4Mux_v I__8087 (
            .O(N__35009),
            .I(N__35002));
    InMux I__8086 (
            .O(N__35008),
            .I(N__34999));
    Span4Mux_v I__8085 (
            .O(N__35005),
            .I(N__34994));
    Span4Mux_h I__8084 (
            .O(N__35002),
            .I(N__34994));
    LocalMux I__8083 (
            .O(N__34999),
            .I(dataRead5_10));
    Odrv4 I__8082 (
            .O(N__34994),
            .I(dataRead5_10));
    InMux I__8081 (
            .O(N__34989),
            .I(N__34986));
    LocalMux I__8080 (
            .O(N__34986),
            .I(N__34983));
    Odrv4 I__8079 (
            .O(N__34983),
            .I(OutReg_0_5_i_m3_ns_1_10));
    CascadeMux I__8078 (
            .O(N__34980),
            .I(N__34975));
    InMux I__8077 (
            .O(N__34979),
            .I(N__34972));
    InMux I__8076 (
            .O(N__34978),
            .I(N__34969));
    InMux I__8075 (
            .O(N__34975),
            .I(N__34966));
    LocalMux I__8074 (
            .O(N__34972),
            .I(N__34961));
    LocalMux I__8073 (
            .O(N__34969),
            .I(N__34961));
    LocalMux I__8072 (
            .O(N__34966),
            .I(N__34958));
    Span4Mux_v I__8071 (
            .O(N__34961),
            .I(N__34953));
    Span4Mux_h I__8070 (
            .O(N__34958),
            .I(N__34953));
    Span4Mux_h I__8069 (
            .O(N__34953),
            .I(N__34950));
    Odrv4 I__8068 (
            .O(N__34950),
            .I(data_receivedZ0Z_4));
    CascadeMux I__8067 (
            .O(N__34947),
            .I(un1_OutReg51_4_0_i_o3_2_cascade_));
    InMux I__8066 (
            .O(N__34944),
            .I(N__34941));
    LocalMux I__8065 (
            .O(N__34941),
            .I(OutReg_21_m_0_a2_1_0));
    InMux I__8064 (
            .O(N__34938),
            .I(N__34935));
    LocalMux I__8063 (
            .O(N__34935),
            .I(OutReg_esr_RNO_2Z0Z_10));
    CascadeMux I__8062 (
            .O(N__34932),
            .I(N__34929));
    InMux I__8061 (
            .O(N__34929),
            .I(N__34926));
    LocalMux I__8060 (
            .O(N__34926),
            .I(N__34923));
    Span4Mux_h I__8059 (
            .O(N__34923),
            .I(N__34920));
    Odrv4 I__8058 (
            .O(N__34920),
            .I(OutRegZ0Z_9));
    InMux I__8057 (
            .O(N__34917),
            .I(N__34914));
    LocalMux I__8056 (
            .O(N__34914),
            .I(OutReg_esr_RNO_0Z0Z_10));
    InMux I__8055 (
            .O(N__34911),
            .I(N__34908));
    LocalMux I__8054 (
            .O(N__34908),
            .I(N__34905));
    Span4Mux_h I__8053 (
            .O(N__34905),
            .I(N__34902));
    Span4Mux_h I__8052 (
            .O(N__34902),
            .I(N__34899));
    Odrv4 I__8051 (
            .O(N__34899),
            .I(OutRegZ0Z_10));
    CascadeMux I__8050 (
            .O(N__34896),
            .I(N__34890));
    InMux I__8049 (
            .O(N__34895),
            .I(N__34886));
    InMux I__8048 (
            .O(N__34894),
            .I(N__34880));
    InMux I__8047 (
            .O(N__34893),
            .I(N__34877));
    InMux I__8046 (
            .O(N__34890),
            .I(N__34874));
    CascadeMux I__8045 (
            .O(N__34889),
            .I(N__34871));
    LocalMux I__8044 (
            .O(N__34886),
            .I(N__34867));
    InMux I__8043 (
            .O(N__34885),
            .I(N__34864));
    CascadeMux I__8042 (
            .O(N__34884),
            .I(N__34859));
    InMux I__8041 (
            .O(N__34883),
            .I(N__34856));
    LocalMux I__8040 (
            .O(N__34880),
            .I(N__34851));
    LocalMux I__8039 (
            .O(N__34877),
            .I(N__34851));
    LocalMux I__8038 (
            .O(N__34874),
            .I(N__34848));
    InMux I__8037 (
            .O(N__34871),
            .I(N__34845));
    InMux I__8036 (
            .O(N__34870),
            .I(N__34842));
    Span4Mux_v I__8035 (
            .O(N__34867),
            .I(N__34839));
    LocalMux I__8034 (
            .O(N__34864),
            .I(N__34836));
    InMux I__8033 (
            .O(N__34863),
            .I(N__34833));
    InMux I__8032 (
            .O(N__34862),
            .I(N__34828));
    InMux I__8031 (
            .O(N__34859),
            .I(N__34828));
    LocalMux I__8030 (
            .O(N__34856),
            .I(N__34823));
    Span4Mux_h I__8029 (
            .O(N__34851),
            .I(N__34823));
    Span4Mux_h I__8028 (
            .O(N__34848),
            .I(N__34818));
    LocalMux I__8027 (
            .O(N__34845),
            .I(N__34818));
    LocalMux I__8026 (
            .O(N__34842),
            .I(data_received_fastZ0Z_2));
    Odrv4 I__8025 (
            .O(N__34839),
            .I(data_received_fastZ0Z_2));
    Odrv12 I__8024 (
            .O(N__34836),
            .I(data_received_fastZ0Z_2));
    LocalMux I__8023 (
            .O(N__34833),
            .I(data_received_fastZ0Z_2));
    LocalMux I__8022 (
            .O(N__34828),
            .I(data_received_fastZ0Z_2));
    Odrv4 I__8021 (
            .O(N__34823),
            .I(data_received_fastZ0Z_2));
    Odrv4 I__8020 (
            .O(N__34818),
            .I(data_received_fastZ0Z_2));
    InMux I__8019 (
            .O(N__34803),
            .I(N__34799));
    InMux I__8018 (
            .O(N__34802),
            .I(N__34796));
    LocalMux I__8017 (
            .O(N__34799),
            .I(N__34793));
    LocalMux I__8016 (
            .O(N__34796),
            .I(N__34790));
    Span4Mux_h I__8015 (
            .O(N__34793),
            .I(N__34784));
    Span4Mux_h I__8014 (
            .O(N__34790),
            .I(N__34784));
    InMux I__8013 (
            .O(N__34789),
            .I(N__34781));
    Span4Mux_h I__8012 (
            .O(N__34784),
            .I(N__34778));
    LocalMux I__8011 (
            .O(N__34781),
            .I(dataRead3_10));
    Odrv4 I__8010 (
            .O(N__34778),
            .I(dataRead3_10));
    CascadeMux I__8009 (
            .O(N__34773),
            .I(N__34768));
    CascadeMux I__8008 (
            .O(N__34772),
            .I(N__34765));
    InMux I__8007 (
            .O(N__34771),
            .I(N__34758));
    InMux I__8006 (
            .O(N__34768),
            .I(N__34755));
    InMux I__8005 (
            .O(N__34765),
            .I(N__34752));
    InMux I__8004 (
            .O(N__34764),
            .I(N__34749));
    InMux I__8003 (
            .O(N__34763),
            .I(N__34746));
    InMux I__8002 (
            .O(N__34762),
            .I(N__34743));
    InMux I__8001 (
            .O(N__34761),
            .I(N__34739));
    LocalMux I__8000 (
            .O(N__34758),
            .I(N__34734));
    LocalMux I__7999 (
            .O(N__34755),
            .I(N__34734));
    LocalMux I__7998 (
            .O(N__34752),
            .I(N__34728));
    LocalMux I__7997 (
            .O(N__34749),
            .I(N__34725));
    LocalMux I__7996 (
            .O(N__34746),
            .I(N__34722));
    LocalMux I__7995 (
            .O(N__34743),
            .I(N__34719));
    InMux I__7994 (
            .O(N__34742),
            .I(N__34716));
    LocalMux I__7993 (
            .O(N__34739),
            .I(N__34711));
    Span4Mux_h I__7992 (
            .O(N__34734),
            .I(N__34711));
    InMux I__7991 (
            .O(N__34733),
            .I(N__34706));
    InMux I__7990 (
            .O(N__34732),
            .I(N__34706));
    InMux I__7989 (
            .O(N__34731),
            .I(N__34703));
    Span4Mux_v I__7988 (
            .O(N__34728),
            .I(N__34696));
    Span4Mux_v I__7987 (
            .O(N__34725),
            .I(N__34696));
    Span4Mux_v I__7986 (
            .O(N__34722),
            .I(N__34696));
    Odrv4 I__7985 (
            .O(N__34719),
            .I(data_received_fastZ0Z_0));
    LocalMux I__7984 (
            .O(N__34716),
            .I(data_received_fastZ0Z_0));
    Odrv4 I__7983 (
            .O(N__34711),
            .I(data_received_fastZ0Z_0));
    LocalMux I__7982 (
            .O(N__34706),
            .I(data_received_fastZ0Z_0));
    LocalMux I__7981 (
            .O(N__34703),
            .I(data_received_fastZ0Z_0));
    Odrv4 I__7980 (
            .O(N__34696),
            .I(data_received_fastZ0Z_0));
    InMux I__7979 (
            .O(N__34683),
            .I(N__34680));
    LocalMux I__7978 (
            .O(N__34680),
            .I(N__34677));
    Span4Mux_v I__7977 (
            .O(N__34677),
            .I(N__34672));
    InMux I__7976 (
            .O(N__34676),
            .I(N__34669));
    InMux I__7975 (
            .O(N__34675),
            .I(N__34666));
    Span4Mux_h I__7974 (
            .O(N__34672),
            .I(N__34663));
    LocalMux I__7973 (
            .O(N__34669),
            .I(N__34660));
    LocalMux I__7972 (
            .O(N__34666),
            .I(N__34655));
    Span4Mux_h I__7971 (
            .O(N__34663),
            .I(N__34655));
    Odrv4 I__7970 (
            .O(N__34660),
            .I(dataRead2_10));
    Odrv4 I__7969 (
            .O(N__34655),
            .I(dataRead2_10));
    InMux I__7968 (
            .O(N__34650),
            .I(N__34646));
    InMux I__7967 (
            .O(N__34649),
            .I(N__34642));
    LocalMux I__7966 (
            .O(N__34646),
            .I(N__34639));
    InMux I__7965 (
            .O(N__34645),
            .I(N__34636));
    LocalMux I__7964 (
            .O(N__34642),
            .I(N__34633));
    Span4Mux_v I__7963 (
            .O(N__34639),
            .I(N__34628));
    LocalMux I__7962 (
            .O(N__34636),
            .I(N__34628));
    Span4Mux_h I__7961 (
            .O(N__34633),
            .I(N__34625));
    Span4Mux_h I__7960 (
            .O(N__34628),
            .I(N__34622));
    Span4Mux_h I__7959 (
            .O(N__34625),
            .I(N__34619));
    Odrv4 I__7958 (
            .O(N__34622),
            .I(dataRead7_10));
    Odrv4 I__7957 (
            .O(N__34619),
            .I(dataRead7_10));
    InMux I__7956 (
            .O(N__34614),
            .I(N__34611));
    LocalMux I__7955 (
            .O(N__34611),
            .I(N__34606));
    InMux I__7954 (
            .O(N__34610),
            .I(N__34603));
    InMux I__7953 (
            .O(N__34609),
            .I(N__34600));
    Span4Mux_h I__7952 (
            .O(N__34606),
            .I(N__34597));
    LocalMux I__7951 (
            .O(N__34603),
            .I(N__34594));
    LocalMux I__7950 (
            .O(N__34600),
            .I(N__34591));
    Span4Mux_h I__7949 (
            .O(N__34597),
            .I(N__34588));
    Odrv4 I__7948 (
            .O(N__34594),
            .I(dataRead6_10));
    Odrv4 I__7947 (
            .O(N__34591),
            .I(dataRead6_10));
    Odrv4 I__7946 (
            .O(N__34588),
            .I(dataRead6_10));
    CascadeMux I__7945 (
            .O(N__34581),
            .I(OutReg_0_4_i_m3_ns_1_10_cascade_));
    InMux I__7944 (
            .O(N__34578),
            .I(N__34575));
    LocalMux I__7943 (
            .O(N__34575),
            .I(OutReg_esr_RNO_1Z0Z_10));
    CascadeMux I__7942 (
            .O(N__34572),
            .I(N__34568));
    InMux I__7941 (
            .O(N__34571),
            .I(N__34564));
    InMux I__7940 (
            .O(N__34568),
            .I(N__34561));
    InMux I__7939 (
            .O(N__34567),
            .I(N__34558));
    LocalMux I__7938 (
            .O(N__34564),
            .I(\PWMInstance2.periodCounter12 ));
    LocalMux I__7937 (
            .O(N__34561),
            .I(\PWMInstance2.periodCounter12 ));
    LocalMux I__7936 (
            .O(N__34558),
            .I(\PWMInstance2.periodCounter12 ));
    InMux I__7935 (
            .O(N__34551),
            .I(N__34546));
    InMux I__7934 (
            .O(N__34550),
            .I(N__34541));
    InMux I__7933 (
            .O(N__34549),
            .I(N__34541));
    LocalMux I__7932 (
            .O(N__34546),
            .I(\PWMInstance2.periodCounterZ0Z_0 ));
    LocalMux I__7931 (
            .O(N__34541),
            .I(\PWMInstance2.periodCounterZ0Z_0 ));
    CascadeMux I__7930 (
            .O(N__34536),
            .I(N__34531));
    CascadeMux I__7929 (
            .O(N__34535),
            .I(N__34528));
    InMux I__7928 (
            .O(N__34534),
            .I(N__34525));
    InMux I__7927 (
            .O(N__34531),
            .I(N__34520));
    InMux I__7926 (
            .O(N__34528),
            .I(N__34520));
    LocalMux I__7925 (
            .O(N__34525),
            .I(\QuadInstance0.delayedCh_AZ0Z_1 ));
    LocalMux I__7924 (
            .O(N__34520),
            .I(\QuadInstance0.delayedCh_AZ0Z_1 ));
    InMux I__7923 (
            .O(N__34515),
            .I(N__34512));
    LocalMux I__7922 (
            .O(N__34512),
            .I(N__34508));
    InMux I__7921 (
            .O(N__34511),
            .I(N__34505));
    Span4Mux_h I__7920 (
            .O(N__34508),
            .I(N__34502));
    LocalMux I__7919 (
            .O(N__34505),
            .I(N__34497));
    Span4Mux_v I__7918 (
            .O(N__34502),
            .I(N__34492));
    InMux I__7917 (
            .O(N__34501),
            .I(N__34489));
    InMux I__7916 (
            .O(N__34500),
            .I(N__34486));
    Span4Mux_v I__7915 (
            .O(N__34497),
            .I(N__34483));
    InMux I__7914 (
            .O(N__34496),
            .I(N__34480));
    InMux I__7913 (
            .O(N__34495),
            .I(N__34477));
    Span4Mux_v I__7912 (
            .O(N__34492),
            .I(N__34472));
    LocalMux I__7911 (
            .O(N__34489),
            .I(N__34472));
    LocalMux I__7910 (
            .O(N__34486),
            .I(N__34466));
    Sp12to4 I__7909 (
            .O(N__34483),
            .I(N__34459));
    LocalMux I__7908 (
            .O(N__34480),
            .I(N__34459));
    LocalMux I__7907 (
            .O(N__34477),
            .I(N__34459));
    Span4Mux_v I__7906 (
            .O(N__34472),
            .I(N__34456));
    InMux I__7905 (
            .O(N__34471),
            .I(N__34453));
    InMux I__7904 (
            .O(N__34470),
            .I(N__34450));
    InMux I__7903 (
            .O(N__34469),
            .I(N__34447));
    Span12Mux_h I__7902 (
            .O(N__34466),
            .I(N__34442));
    Span12Mux_h I__7901 (
            .O(N__34459),
            .I(N__34442));
    Span4Mux_v I__7900 (
            .O(N__34456),
            .I(N__34439));
    LocalMux I__7899 (
            .O(N__34453),
            .I(N__34432));
    LocalMux I__7898 (
            .O(N__34450),
            .I(N__34432));
    LocalMux I__7897 (
            .O(N__34447),
            .I(N__34432));
    Span12Mux_v I__7896 (
            .O(N__34442),
            .I(N__34429));
    IoSpan4Mux I__7895 (
            .O(N__34439),
            .I(N__34426));
    Span12Mux_h I__7894 (
            .O(N__34432),
            .I(N__34423));
    Odrv12 I__7893 (
            .O(N__34429),
            .I(RST_c));
    Odrv4 I__7892 (
            .O(N__34426),
            .I(RST_c));
    Odrv12 I__7891 (
            .O(N__34423),
            .I(RST_c));
    InMux I__7890 (
            .O(N__34416),
            .I(N__34410));
    InMux I__7889 (
            .O(N__34415),
            .I(N__34407));
    InMux I__7888 (
            .O(N__34414),
            .I(N__34404));
    InMux I__7887 (
            .O(N__34413),
            .I(N__34396));
    LocalMux I__7886 (
            .O(N__34410),
            .I(N__34391));
    LocalMux I__7885 (
            .O(N__34407),
            .I(N__34388));
    LocalMux I__7884 (
            .O(N__34404),
            .I(N__34385));
    InMux I__7883 (
            .O(N__34403),
            .I(N__34382));
    InMux I__7882 (
            .O(N__34402),
            .I(N__34379));
    InMux I__7881 (
            .O(N__34401),
            .I(N__34375));
    InMux I__7880 (
            .O(N__34400),
            .I(N__34370));
    InMux I__7879 (
            .O(N__34399),
            .I(N__34367));
    LocalMux I__7878 (
            .O(N__34396),
            .I(N__34362));
    InMux I__7877 (
            .O(N__34395),
            .I(N__34359));
    InMux I__7876 (
            .O(N__34394),
            .I(N__34356));
    Span4Mux_v I__7875 (
            .O(N__34391),
            .I(N__34351));
    Span4Mux_h I__7874 (
            .O(N__34388),
            .I(N__34351));
    Span4Mux_h I__7873 (
            .O(N__34385),
            .I(N__34346));
    LocalMux I__7872 (
            .O(N__34382),
            .I(N__34346));
    LocalMux I__7871 (
            .O(N__34379),
            .I(N__34343));
    InMux I__7870 (
            .O(N__34378),
            .I(N__34340));
    LocalMux I__7869 (
            .O(N__34375),
            .I(N__34337));
    InMux I__7868 (
            .O(N__34374),
            .I(N__34332));
    InMux I__7867 (
            .O(N__34373),
            .I(N__34332));
    LocalMux I__7866 (
            .O(N__34370),
            .I(N__34329));
    LocalMux I__7865 (
            .O(N__34367),
            .I(N__34326));
    InMux I__7864 (
            .O(N__34366),
            .I(N__34323));
    InMux I__7863 (
            .O(N__34365),
            .I(N__34320));
    Span4Mux_v I__7862 (
            .O(N__34362),
            .I(N__34317));
    LocalMux I__7861 (
            .O(N__34359),
            .I(N__34312));
    LocalMux I__7860 (
            .O(N__34356),
            .I(N__34312));
    Span4Mux_v I__7859 (
            .O(N__34351),
            .I(N__34309));
    Span4Mux_h I__7858 (
            .O(N__34346),
            .I(N__34304));
    Span4Mux_h I__7857 (
            .O(N__34343),
            .I(N__34304));
    LocalMux I__7856 (
            .O(N__34340),
            .I(N__34301));
    Span4Mux_v I__7855 (
            .O(N__34337),
            .I(N__34298));
    LocalMux I__7854 (
            .O(N__34332),
            .I(N__34295));
    Span4Mux_h I__7853 (
            .O(N__34329),
            .I(N__34292));
    Span4Mux_h I__7852 (
            .O(N__34326),
            .I(N__34285));
    LocalMux I__7851 (
            .O(N__34323),
            .I(N__34285));
    LocalMux I__7850 (
            .O(N__34320),
            .I(N__34285));
    Span4Mux_h I__7849 (
            .O(N__34317),
            .I(N__34276));
    Span4Mux_v I__7848 (
            .O(N__34312),
            .I(N__34276));
    Span4Mux_h I__7847 (
            .O(N__34309),
            .I(N__34276));
    Span4Mux_v I__7846 (
            .O(N__34304),
            .I(N__34276));
    Span4Mux_h I__7845 (
            .O(N__34301),
            .I(N__34269));
    Span4Mux_h I__7844 (
            .O(N__34298),
            .I(N__34269));
    Span4Mux_v I__7843 (
            .O(N__34295),
            .I(N__34269));
    Span4Mux_h I__7842 (
            .O(N__34292),
            .I(N__34264));
    Span4Mux_h I__7841 (
            .O(N__34285),
            .I(N__34264));
    Odrv4 I__7840 (
            .O(N__34276),
            .I(dataWriteZ0Z_14));
    Odrv4 I__7839 (
            .O(N__34269),
            .I(dataWriteZ0Z_14));
    Odrv4 I__7838 (
            .O(N__34264),
            .I(dataWriteZ0Z_14));
    InMux I__7837 (
            .O(N__34257),
            .I(N__34254));
    LocalMux I__7836 (
            .O(N__34254),
            .I(\QuadInstance0.Quad_RNO_0_0_14 ));
    InMux I__7835 (
            .O(N__34251),
            .I(N__34246));
    CascadeMux I__7834 (
            .O(N__34250),
            .I(N__34243));
    InMux I__7833 (
            .O(N__34249),
            .I(N__34240));
    LocalMux I__7832 (
            .O(N__34246),
            .I(N__34237));
    InMux I__7831 (
            .O(N__34243),
            .I(N__34234));
    LocalMux I__7830 (
            .O(N__34240),
            .I(N__34229));
    Span4Mux_v I__7829 (
            .O(N__34237),
            .I(N__34229));
    LocalMux I__7828 (
            .O(N__34234),
            .I(dataRead0_14));
    Odrv4 I__7827 (
            .O(N__34229),
            .I(dataRead0_14));
    InMux I__7826 (
            .O(N__34224),
            .I(N__34221));
    LocalMux I__7825 (
            .O(N__34221),
            .I(\QuadInstance0.Quad_RNI4P8Q1Z0Z_14 ));
    CascadeMux I__7824 (
            .O(N__34218),
            .I(N__34214));
    InMux I__7823 (
            .O(N__34217),
            .I(N__34211));
    InMux I__7822 (
            .O(N__34214),
            .I(N__34208));
    LocalMux I__7821 (
            .O(N__34211),
            .I(N__34204));
    LocalMux I__7820 (
            .O(N__34208),
            .I(N__34201));
    InMux I__7819 (
            .O(N__34207),
            .I(N__34198));
    Span4Mux_h I__7818 (
            .O(N__34204),
            .I(N__34195));
    Span4Mux_h I__7817 (
            .O(N__34201),
            .I(N__34192));
    LocalMux I__7816 (
            .O(N__34198),
            .I(N__34189));
    Span4Mux_h I__7815 (
            .O(N__34195),
            .I(N__34186));
    Span4Mux_h I__7814 (
            .O(N__34192),
            .I(N__34183));
    Odrv12 I__7813 (
            .O(N__34189),
            .I(dataRead0_3));
    Odrv4 I__7812 (
            .O(N__34186),
            .I(dataRead0_3));
    Odrv4 I__7811 (
            .O(N__34183),
            .I(dataRead0_3));
    InMux I__7810 (
            .O(N__34176),
            .I(N__34173));
    LocalMux I__7809 (
            .O(N__34173),
            .I(\QuadInstance0.Quad_RNIIGBH1Z0Z_3 ));
    CascadeMux I__7808 (
            .O(N__34170),
            .I(N__34167));
    InMux I__7807 (
            .O(N__34167),
            .I(N__34164));
    LocalMux I__7806 (
            .O(N__34164),
            .I(N__34160));
    InMux I__7805 (
            .O(N__34163),
            .I(N__34157));
    Span4Mux_v I__7804 (
            .O(N__34160),
            .I(N__34154));
    LocalMux I__7803 (
            .O(N__34157),
            .I(N__34150));
    Sp12to4 I__7802 (
            .O(N__34154),
            .I(N__34147));
    InMux I__7801 (
            .O(N__34153),
            .I(N__34144));
    Span4Mux_v I__7800 (
            .O(N__34150),
            .I(N__34141));
    Odrv12 I__7799 (
            .O(N__34147),
            .I(dataRead0_4));
    LocalMux I__7798 (
            .O(N__34144),
            .I(dataRead0_4));
    Odrv4 I__7797 (
            .O(N__34141),
            .I(dataRead0_4));
    CascadeMux I__7796 (
            .O(N__34134),
            .I(N__34131));
    InMux I__7795 (
            .O(N__34131),
            .I(N__34128));
    LocalMux I__7794 (
            .O(N__34128),
            .I(\QuadInstance0.Quad_RNIJHBH1Z0Z_4 ));
    InMux I__7793 (
            .O(N__34125),
            .I(N__34122));
    LocalMux I__7792 (
            .O(N__34122),
            .I(N__34118));
    InMux I__7791 (
            .O(N__34121),
            .I(N__34115));
    Span4Mux_v I__7790 (
            .O(N__34118),
            .I(N__34111));
    LocalMux I__7789 (
            .O(N__34115),
            .I(N__34108));
    InMux I__7788 (
            .O(N__34114),
            .I(N__34105));
    Odrv4 I__7787 (
            .O(N__34111),
            .I(dataRead0_5));
    Odrv4 I__7786 (
            .O(N__34108),
            .I(dataRead0_5));
    LocalMux I__7785 (
            .O(N__34105),
            .I(dataRead0_5));
    CascadeMux I__7784 (
            .O(N__34098),
            .I(N__34095));
    InMux I__7783 (
            .O(N__34095),
            .I(N__34092));
    LocalMux I__7782 (
            .O(N__34092),
            .I(\QuadInstance0.Quad_RNIKIBH1Z0Z_5 ));
    InMux I__7781 (
            .O(N__34089),
            .I(N__34082));
    CascadeMux I__7780 (
            .O(N__34088),
            .I(N__34078));
    CascadeMux I__7779 (
            .O(N__34087),
            .I(N__34074));
    CascadeMux I__7778 (
            .O(N__34086),
            .I(N__34071));
    CascadeMux I__7777 (
            .O(N__34085),
            .I(N__34068));
    LocalMux I__7776 (
            .O(N__34082),
            .I(N__34065));
    CascadeMux I__7775 (
            .O(N__34081),
            .I(N__34062));
    InMux I__7774 (
            .O(N__34078),
            .I(N__34054));
    InMux I__7773 (
            .O(N__34077),
            .I(N__34054));
    InMux I__7772 (
            .O(N__34074),
            .I(N__34054));
    InMux I__7771 (
            .O(N__34071),
            .I(N__34049));
    InMux I__7770 (
            .O(N__34068),
            .I(N__34049));
    Span4Mux_v I__7769 (
            .O(N__34065),
            .I(N__34043));
    InMux I__7768 (
            .O(N__34062),
            .I(N__34038));
    InMux I__7767 (
            .O(N__34061),
            .I(N__34038));
    LocalMux I__7766 (
            .O(N__34054),
            .I(N__34033));
    LocalMux I__7765 (
            .O(N__34049),
            .I(N__34033));
    CascadeMux I__7764 (
            .O(N__34048),
            .I(N__34025));
    InMux I__7763 (
            .O(N__34047),
            .I(N__34022));
    InMux I__7762 (
            .O(N__34046),
            .I(N__34019));
    Span4Mux_h I__7761 (
            .O(N__34043),
            .I(N__34014));
    LocalMux I__7760 (
            .O(N__34038),
            .I(N__34014));
    Span4Mux_h I__7759 (
            .O(N__34033),
            .I(N__34011));
    InMux I__7758 (
            .O(N__34032),
            .I(N__34002));
    InMux I__7757 (
            .O(N__34031),
            .I(N__34002));
    InMux I__7756 (
            .O(N__34030),
            .I(N__34002));
    InMux I__7755 (
            .O(N__34029),
            .I(N__34002));
    InMux I__7754 (
            .O(N__34028),
            .I(N__33997));
    InMux I__7753 (
            .O(N__34025),
            .I(N__33997));
    LocalMux I__7752 (
            .O(N__34022),
            .I(\QuadInstance0.count_enable ));
    LocalMux I__7751 (
            .O(N__34019),
            .I(\QuadInstance0.count_enable ));
    Odrv4 I__7750 (
            .O(N__34014),
            .I(\QuadInstance0.count_enable ));
    Odrv4 I__7749 (
            .O(N__34011),
            .I(\QuadInstance0.count_enable ));
    LocalMux I__7748 (
            .O(N__34002),
            .I(\QuadInstance0.count_enable ));
    LocalMux I__7747 (
            .O(N__33997),
            .I(\QuadInstance0.count_enable ));
    CascadeMux I__7746 (
            .O(N__33984),
            .I(N__33981));
    InMux I__7745 (
            .O(N__33981),
            .I(N__33977));
    InMux I__7744 (
            .O(N__33980),
            .I(N__33974));
    LocalMux I__7743 (
            .O(N__33977),
            .I(N__33971));
    LocalMux I__7742 (
            .O(N__33974),
            .I(N__33967));
    Span4Mux_v I__7741 (
            .O(N__33971),
            .I(N__33964));
    InMux I__7740 (
            .O(N__33970),
            .I(N__33961));
    Span4Mux_h I__7739 (
            .O(N__33967),
            .I(N__33958));
    Odrv4 I__7738 (
            .O(N__33964),
            .I(dataRead0_6));
    LocalMux I__7737 (
            .O(N__33961),
            .I(dataRead0_6));
    Odrv4 I__7736 (
            .O(N__33958),
            .I(dataRead0_6));
    CascadeMux I__7735 (
            .O(N__33951),
            .I(N__33946));
    CascadeMux I__7734 (
            .O(N__33950),
            .I(N__33939));
    InMux I__7733 (
            .O(N__33949),
            .I(N__33932));
    InMux I__7732 (
            .O(N__33946),
            .I(N__33932));
    InMux I__7731 (
            .O(N__33945),
            .I(N__33932));
    InMux I__7730 (
            .O(N__33944),
            .I(N__33927));
    InMux I__7729 (
            .O(N__33943),
            .I(N__33927));
    InMux I__7728 (
            .O(N__33942),
            .I(N__33919));
    InMux I__7727 (
            .O(N__33939),
            .I(N__33919));
    LocalMux I__7726 (
            .O(N__33932),
            .I(N__33914));
    LocalMux I__7725 (
            .O(N__33927),
            .I(N__33914));
    CascadeMux I__7724 (
            .O(N__33926),
            .I(N__33910));
    CascadeMux I__7723 (
            .O(N__33925),
            .I(N__33906));
    InMux I__7722 (
            .O(N__33924),
            .I(N__33900));
    LocalMux I__7721 (
            .O(N__33919),
            .I(N__33897));
    Span4Mux_h I__7720 (
            .O(N__33914),
            .I(N__33894));
    InMux I__7719 (
            .O(N__33913),
            .I(N__33883));
    InMux I__7718 (
            .O(N__33910),
            .I(N__33883));
    InMux I__7717 (
            .O(N__33909),
            .I(N__33883));
    InMux I__7716 (
            .O(N__33906),
            .I(N__33883));
    InMux I__7715 (
            .O(N__33905),
            .I(N__33883));
    InMux I__7714 (
            .O(N__33904),
            .I(N__33878));
    InMux I__7713 (
            .O(N__33903),
            .I(N__33878));
    LocalMux I__7712 (
            .O(N__33900),
            .I(\QuadInstance0.un1_count_enable_i_a2_0_1 ));
    Odrv4 I__7711 (
            .O(N__33897),
            .I(\QuadInstance0.un1_count_enable_i_a2_0_1 ));
    Odrv4 I__7710 (
            .O(N__33894),
            .I(\QuadInstance0.un1_count_enable_i_a2_0_1 ));
    LocalMux I__7709 (
            .O(N__33883),
            .I(\QuadInstance0.un1_count_enable_i_a2_0_1 ));
    LocalMux I__7708 (
            .O(N__33878),
            .I(\QuadInstance0.un1_count_enable_i_a2_0_1 ));
    CascadeMux I__7707 (
            .O(N__33867),
            .I(N__33864));
    InMux I__7706 (
            .O(N__33864),
            .I(N__33861));
    LocalMux I__7705 (
            .O(N__33861),
            .I(\QuadInstance0.Quad_RNILJBH1Z0Z_6 ));
    InMux I__7704 (
            .O(N__33858),
            .I(N__33852));
    InMux I__7703 (
            .O(N__33857),
            .I(N__33843));
    InMux I__7702 (
            .O(N__33856),
            .I(N__33837));
    InMux I__7701 (
            .O(N__33855),
            .I(N__33837));
    LocalMux I__7700 (
            .O(N__33852),
            .I(N__33834));
    InMux I__7699 (
            .O(N__33851),
            .I(N__33831));
    InMux I__7698 (
            .O(N__33850),
            .I(N__33823));
    InMux I__7697 (
            .O(N__33849),
            .I(N__33819));
    InMux I__7696 (
            .O(N__33848),
            .I(N__33816));
    InMux I__7695 (
            .O(N__33847),
            .I(N__33813));
    InMux I__7694 (
            .O(N__33846),
            .I(N__33810));
    LocalMux I__7693 (
            .O(N__33843),
            .I(N__33807));
    InMux I__7692 (
            .O(N__33842),
            .I(N__33804));
    LocalMux I__7691 (
            .O(N__33837),
            .I(N__33801));
    Span4Mux_v I__7690 (
            .O(N__33834),
            .I(N__33796));
    LocalMux I__7689 (
            .O(N__33831),
            .I(N__33796));
    InMux I__7688 (
            .O(N__33830),
            .I(N__33793));
    InMux I__7687 (
            .O(N__33829),
            .I(N__33788));
    InMux I__7686 (
            .O(N__33828),
            .I(N__33788));
    InMux I__7685 (
            .O(N__33827),
            .I(N__33785));
    InMux I__7684 (
            .O(N__33826),
            .I(N__33780));
    LocalMux I__7683 (
            .O(N__33823),
            .I(N__33777));
    InMux I__7682 (
            .O(N__33822),
            .I(N__33774));
    LocalMux I__7681 (
            .O(N__33819),
            .I(N__33771));
    LocalMux I__7680 (
            .O(N__33816),
            .I(N__33762));
    LocalMux I__7679 (
            .O(N__33813),
            .I(N__33762));
    LocalMux I__7678 (
            .O(N__33810),
            .I(N__33762));
    Span4Mux_h I__7677 (
            .O(N__33807),
            .I(N__33762));
    LocalMux I__7676 (
            .O(N__33804),
            .I(N__33752));
    Span4Mux_v I__7675 (
            .O(N__33801),
            .I(N__33752));
    Span4Mux_h I__7674 (
            .O(N__33796),
            .I(N__33752));
    LocalMux I__7673 (
            .O(N__33793),
            .I(N__33744));
    LocalMux I__7672 (
            .O(N__33788),
            .I(N__33744));
    LocalMux I__7671 (
            .O(N__33785),
            .I(N__33741));
    InMux I__7670 (
            .O(N__33784),
            .I(N__33736));
    InMux I__7669 (
            .O(N__33783),
            .I(N__33736));
    LocalMux I__7668 (
            .O(N__33780),
            .I(N__33733));
    Span4Mux_v I__7667 (
            .O(N__33777),
            .I(N__33730));
    LocalMux I__7666 (
            .O(N__33774),
            .I(N__33723));
    Span4Mux_v I__7665 (
            .O(N__33771),
            .I(N__33723));
    Span4Mux_v I__7664 (
            .O(N__33762),
            .I(N__33723));
    InMux I__7663 (
            .O(N__33761),
            .I(N__33716));
    InMux I__7662 (
            .O(N__33760),
            .I(N__33716));
    InMux I__7661 (
            .O(N__33759),
            .I(N__33716));
    Span4Mux_v I__7660 (
            .O(N__33752),
            .I(N__33713));
    InMux I__7659 (
            .O(N__33751),
            .I(N__33708));
    InMux I__7658 (
            .O(N__33750),
            .I(N__33708));
    InMux I__7657 (
            .O(N__33749),
            .I(N__33705));
    Span4Mux_h I__7656 (
            .O(N__33744),
            .I(N__33702));
    Span12Mux_s11_v I__7655 (
            .O(N__33741),
            .I(N__33699));
    LocalMux I__7654 (
            .O(N__33736),
            .I(N__33690));
    Span4Mux_v I__7653 (
            .O(N__33733),
            .I(N__33690));
    Span4Mux_h I__7652 (
            .O(N__33730),
            .I(N__33690));
    Span4Mux_h I__7651 (
            .O(N__33723),
            .I(N__33690));
    LocalMux I__7650 (
            .O(N__33716),
            .I(N__33685));
    Span4Mux_h I__7649 (
            .O(N__33713),
            .I(N__33685));
    LocalMux I__7648 (
            .O(N__33708),
            .I(data_receivedZ0Z_21));
    LocalMux I__7647 (
            .O(N__33705),
            .I(data_receivedZ0Z_21));
    Odrv4 I__7646 (
            .O(N__33702),
            .I(data_receivedZ0Z_21));
    Odrv12 I__7645 (
            .O(N__33699),
            .I(data_receivedZ0Z_21));
    Odrv4 I__7644 (
            .O(N__33690),
            .I(data_receivedZ0Z_21));
    Odrv4 I__7643 (
            .O(N__33685),
            .I(data_receivedZ0Z_21));
    InMux I__7642 (
            .O(N__33672),
            .I(N__33667));
    CascadeMux I__7641 (
            .O(N__33671),
            .I(N__33663));
    InMux I__7640 (
            .O(N__33670),
            .I(N__33653));
    LocalMux I__7639 (
            .O(N__33667),
            .I(N__33648));
    InMux I__7638 (
            .O(N__33666),
            .I(N__33645));
    InMux I__7637 (
            .O(N__33663),
            .I(N__33640));
    InMux I__7636 (
            .O(N__33662),
            .I(N__33640));
    CascadeMux I__7635 (
            .O(N__33661),
            .I(N__33634));
    InMux I__7634 (
            .O(N__33660),
            .I(N__33631));
    InMux I__7633 (
            .O(N__33659),
            .I(N__33628));
    InMux I__7632 (
            .O(N__33658),
            .I(N__33623));
    InMux I__7631 (
            .O(N__33657),
            .I(N__33623));
    InMux I__7630 (
            .O(N__33656),
            .I(N__33620));
    LocalMux I__7629 (
            .O(N__33653),
            .I(N__33616));
    InMux I__7628 (
            .O(N__33652),
            .I(N__33611));
    InMux I__7627 (
            .O(N__33651),
            .I(N__33611));
    Span4Mux_v I__7626 (
            .O(N__33648),
            .I(N__33604));
    LocalMux I__7625 (
            .O(N__33645),
            .I(N__33604));
    LocalMux I__7624 (
            .O(N__33640),
            .I(N__33604));
    InMux I__7623 (
            .O(N__33639),
            .I(N__33601));
    CascadeMux I__7622 (
            .O(N__33638),
            .I(N__33596));
    CascadeMux I__7621 (
            .O(N__33637),
            .I(N__33593));
    InMux I__7620 (
            .O(N__33634),
            .I(N__33590));
    LocalMux I__7619 (
            .O(N__33631),
            .I(N__33587));
    LocalMux I__7618 (
            .O(N__33628),
            .I(N__33583));
    LocalMux I__7617 (
            .O(N__33623),
            .I(N__33578));
    LocalMux I__7616 (
            .O(N__33620),
            .I(N__33578));
    InMux I__7615 (
            .O(N__33619),
            .I(N__33575));
    Span4Mux_v I__7614 (
            .O(N__33616),
            .I(N__33572));
    LocalMux I__7613 (
            .O(N__33611),
            .I(N__33565));
    Span4Mux_v I__7612 (
            .O(N__33604),
            .I(N__33565));
    LocalMux I__7611 (
            .O(N__33601),
            .I(N__33565));
    CascadeMux I__7610 (
            .O(N__33600),
            .I(N__33562));
    InMux I__7609 (
            .O(N__33599),
            .I(N__33554));
    InMux I__7608 (
            .O(N__33596),
            .I(N__33549));
    InMux I__7607 (
            .O(N__33593),
            .I(N__33549));
    LocalMux I__7606 (
            .O(N__33590),
            .I(N__33546));
    Span4Mux_v I__7605 (
            .O(N__33587),
            .I(N__33543));
    InMux I__7604 (
            .O(N__33586),
            .I(N__33540));
    Span4Mux_v I__7603 (
            .O(N__33583),
            .I(N__33537));
    Span4Mux_v I__7602 (
            .O(N__33578),
            .I(N__33534));
    LocalMux I__7601 (
            .O(N__33575),
            .I(N__33531));
    Span4Mux_h I__7600 (
            .O(N__33572),
            .I(N__33526));
    Span4Mux_v I__7599 (
            .O(N__33565),
            .I(N__33526));
    InMux I__7598 (
            .O(N__33562),
            .I(N__33521));
    InMux I__7597 (
            .O(N__33561),
            .I(N__33521));
    InMux I__7596 (
            .O(N__33560),
            .I(N__33518));
    InMux I__7595 (
            .O(N__33559),
            .I(N__33511));
    InMux I__7594 (
            .O(N__33558),
            .I(N__33511));
    InMux I__7593 (
            .O(N__33557),
            .I(N__33511));
    LocalMux I__7592 (
            .O(N__33554),
            .I(N__33508));
    LocalMux I__7591 (
            .O(N__33549),
            .I(N__33503));
    Span4Mux_h I__7590 (
            .O(N__33546),
            .I(N__33503));
    Span4Mux_h I__7589 (
            .O(N__33543),
            .I(N__33500));
    LocalMux I__7588 (
            .O(N__33540),
            .I(N__33493));
    Span4Mux_h I__7587 (
            .O(N__33537),
            .I(N__33493));
    Span4Mux_v I__7586 (
            .O(N__33534),
            .I(N__33493));
    Span12Mux_s11_v I__7585 (
            .O(N__33531),
            .I(N__33490));
    Span4Mux_h I__7584 (
            .O(N__33526),
            .I(N__33487));
    LocalMux I__7583 (
            .O(N__33521),
            .I(data_receivedZ0Z_20));
    LocalMux I__7582 (
            .O(N__33518),
            .I(data_receivedZ0Z_20));
    LocalMux I__7581 (
            .O(N__33511),
            .I(data_receivedZ0Z_20));
    Odrv4 I__7580 (
            .O(N__33508),
            .I(data_receivedZ0Z_20));
    Odrv4 I__7579 (
            .O(N__33503),
            .I(data_receivedZ0Z_20));
    Odrv4 I__7578 (
            .O(N__33500),
            .I(data_receivedZ0Z_20));
    Odrv4 I__7577 (
            .O(N__33493),
            .I(data_receivedZ0Z_20));
    Odrv12 I__7576 (
            .O(N__33490),
            .I(data_receivedZ0Z_20));
    Odrv4 I__7575 (
            .O(N__33487),
            .I(data_receivedZ0Z_20));
    CascadeMux I__7574 (
            .O(N__33468),
            .I(N__33460));
    CascadeMux I__7573 (
            .O(N__33467),
            .I(N__33453));
    CascadeMux I__7572 (
            .O(N__33466),
            .I(N__33443));
    CascadeMux I__7571 (
            .O(N__33465),
            .I(N__33437));
    CascadeMux I__7570 (
            .O(N__33464),
            .I(N__33433));
    CascadeMux I__7569 (
            .O(N__33463),
            .I(N__33429));
    InMux I__7568 (
            .O(N__33460),
            .I(N__33426));
    InMux I__7567 (
            .O(N__33459),
            .I(N__33421));
    InMux I__7566 (
            .O(N__33458),
            .I(N__33421));
    InMux I__7565 (
            .O(N__33457),
            .I(N__33416));
    InMux I__7564 (
            .O(N__33456),
            .I(N__33416));
    InMux I__7563 (
            .O(N__33453),
            .I(N__33413));
    CascadeMux I__7562 (
            .O(N__33452),
            .I(N__33410));
    CascadeMux I__7561 (
            .O(N__33451),
            .I(N__33407));
    CascadeMux I__7560 (
            .O(N__33450),
            .I(N__33404));
    CascadeMux I__7559 (
            .O(N__33449),
            .I(N__33401));
    CascadeMux I__7558 (
            .O(N__33448),
            .I(N__33397));
    CascadeMux I__7557 (
            .O(N__33447),
            .I(N__33394));
    CascadeMux I__7556 (
            .O(N__33446),
            .I(N__33391));
    InMux I__7555 (
            .O(N__33443),
            .I(N__33388));
    CascadeMux I__7554 (
            .O(N__33442),
            .I(N__33385));
    CascadeMux I__7553 (
            .O(N__33441),
            .I(N__33382));
    InMux I__7552 (
            .O(N__33440),
            .I(N__33377));
    InMux I__7551 (
            .O(N__33437),
            .I(N__33377));
    InMux I__7550 (
            .O(N__33436),
            .I(N__33374));
    InMux I__7549 (
            .O(N__33433),
            .I(N__33371));
    CascadeMux I__7548 (
            .O(N__33432),
            .I(N__33368));
    InMux I__7547 (
            .O(N__33429),
            .I(N__33364));
    LocalMux I__7546 (
            .O(N__33426),
            .I(N__33357));
    LocalMux I__7545 (
            .O(N__33421),
            .I(N__33357));
    LocalMux I__7544 (
            .O(N__33416),
            .I(N__33357));
    LocalMux I__7543 (
            .O(N__33413),
            .I(N__33354));
    InMux I__7542 (
            .O(N__33410),
            .I(N__33351));
    InMux I__7541 (
            .O(N__33407),
            .I(N__33346));
    InMux I__7540 (
            .O(N__33404),
            .I(N__33346));
    InMux I__7539 (
            .O(N__33401),
            .I(N__33343));
    CascadeMux I__7538 (
            .O(N__33400),
            .I(N__33340));
    InMux I__7537 (
            .O(N__33397),
            .I(N__33337));
    InMux I__7536 (
            .O(N__33394),
            .I(N__33332));
    InMux I__7535 (
            .O(N__33391),
            .I(N__33332));
    LocalMux I__7534 (
            .O(N__33388),
            .I(N__33329));
    InMux I__7533 (
            .O(N__33385),
            .I(N__33326));
    InMux I__7532 (
            .O(N__33382),
            .I(N__33323));
    LocalMux I__7531 (
            .O(N__33377),
            .I(N__33316));
    LocalMux I__7530 (
            .O(N__33374),
            .I(N__33316));
    LocalMux I__7529 (
            .O(N__33371),
            .I(N__33316));
    InMux I__7528 (
            .O(N__33368),
            .I(N__33311));
    InMux I__7527 (
            .O(N__33367),
            .I(N__33311));
    LocalMux I__7526 (
            .O(N__33364),
            .I(N__33304));
    Span4Mux_v I__7525 (
            .O(N__33357),
            .I(N__33304));
    Span4Mux_v I__7524 (
            .O(N__33354),
            .I(N__33304));
    LocalMux I__7523 (
            .O(N__33351),
            .I(N__33301));
    LocalMux I__7522 (
            .O(N__33346),
            .I(N__33298));
    LocalMux I__7521 (
            .O(N__33343),
            .I(N__33295));
    InMux I__7520 (
            .O(N__33340),
            .I(N__33292));
    LocalMux I__7519 (
            .O(N__33337),
            .I(N__33287));
    LocalMux I__7518 (
            .O(N__33332),
            .I(N__33287));
    Span4Mux_h I__7517 (
            .O(N__33329),
            .I(N__33284));
    LocalMux I__7516 (
            .O(N__33326),
            .I(N__33276));
    LocalMux I__7515 (
            .O(N__33323),
            .I(N__33276));
    Span4Mux_v I__7514 (
            .O(N__33316),
            .I(N__33276));
    LocalMux I__7513 (
            .O(N__33311),
            .I(N__33267));
    Span4Mux_h I__7512 (
            .O(N__33304),
            .I(N__33267));
    Span4Mux_v I__7511 (
            .O(N__33301),
            .I(N__33267));
    Span4Mux_v I__7510 (
            .O(N__33298),
            .I(N__33267));
    Sp12to4 I__7509 (
            .O(N__33295),
            .I(N__33264));
    LocalMux I__7508 (
            .O(N__33292),
            .I(N__33259));
    Span4Mux_h I__7507 (
            .O(N__33287),
            .I(N__33259));
    Span4Mux_v I__7506 (
            .O(N__33284),
            .I(N__33256));
    InMux I__7505 (
            .O(N__33283),
            .I(N__33253));
    Sp12to4 I__7504 (
            .O(N__33276),
            .I(N__33246));
    Sp12to4 I__7503 (
            .O(N__33267),
            .I(N__33246));
    Span12Mux_s9_v I__7502 (
            .O(N__33264),
            .I(N__33246));
    Span4Mux_v I__7501 (
            .O(N__33259),
            .I(N__33241));
    Span4Mux_h I__7500 (
            .O(N__33256),
            .I(N__33241));
    LocalMux I__7499 (
            .O(N__33253),
            .I(data_receivedZ0Z_22));
    Odrv12 I__7498 (
            .O(N__33246),
            .I(data_receivedZ0Z_22));
    Odrv4 I__7497 (
            .O(N__33241),
            .I(data_receivedZ0Z_22));
    InMux I__7496 (
            .O(N__33234),
            .I(N__33226));
    InMux I__7495 (
            .O(N__33233),
            .I(N__33226));
    InMux I__7494 (
            .O(N__33232),
            .I(N__33221));
    InMux I__7493 (
            .O(N__33231),
            .I(N__33218));
    LocalMux I__7492 (
            .O(N__33226),
            .I(N__33215));
    InMux I__7491 (
            .O(N__33225),
            .I(N__33211));
    InMux I__7490 (
            .O(N__33224),
            .I(N__33208));
    LocalMux I__7489 (
            .O(N__33221),
            .I(N__33204));
    LocalMux I__7488 (
            .O(N__33218),
            .I(N__33200));
    Span4Mux_h I__7487 (
            .O(N__33215),
            .I(N__33197));
    InMux I__7486 (
            .O(N__33214),
            .I(N__33194));
    LocalMux I__7485 (
            .O(N__33211),
            .I(N__33189));
    LocalMux I__7484 (
            .O(N__33208),
            .I(N__33186));
    InMux I__7483 (
            .O(N__33207),
            .I(N__33183));
    Span4Mux_h I__7482 (
            .O(N__33204),
            .I(N__33180));
    InMux I__7481 (
            .O(N__33203),
            .I(N__33177));
    Span4Mux_h I__7480 (
            .O(N__33200),
            .I(N__33174));
    Span4Mux_v I__7479 (
            .O(N__33197),
            .I(N__33169));
    LocalMux I__7478 (
            .O(N__33194),
            .I(N__33169));
    InMux I__7477 (
            .O(N__33193),
            .I(N__33164));
    InMux I__7476 (
            .O(N__33192),
            .I(N__33164));
    Span4Mux_v I__7475 (
            .O(N__33189),
            .I(N__33157));
    Span4Mux_v I__7474 (
            .O(N__33186),
            .I(N__33157));
    LocalMux I__7473 (
            .O(N__33183),
            .I(N__33157));
    Span4Mux_h I__7472 (
            .O(N__33180),
            .I(N__33154));
    LocalMux I__7471 (
            .O(N__33177),
            .I(N__33151));
    Span4Mux_h I__7470 (
            .O(N__33174),
            .I(N__33144));
    Span4Mux_h I__7469 (
            .O(N__33169),
            .I(N__33144));
    LocalMux I__7468 (
            .O(N__33164),
            .I(N__33144));
    Span4Mux_h I__7467 (
            .O(N__33157),
            .I(N__33141));
    Odrv4 I__7466 (
            .O(N__33154),
            .I(data_received_esr_RNIMIH31_0Z0Z_19));
    Odrv4 I__7465 (
            .O(N__33151),
            .I(data_received_esr_RNIMIH31_0Z0Z_19));
    Odrv4 I__7464 (
            .O(N__33144),
            .I(data_received_esr_RNIMIH31_0Z0Z_19));
    Odrv4 I__7463 (
            .O(N__33141),
            .I(data_received_esr_RNIMIH31_0Z0Z_19));
    InMux I__7462 (
            .O(N__33132),
            .I(N__33121));
    InMux I__7461 (
            .O(N__33131),
            .I(N__33121));
    InMux I__7460 (
            .O(N__33130),
            .I(N__33117));
    InMux I__7459 (
            .O(N__33129),
            .I(N__33104));
    InMux I__7458 (
            .O(N__33128),
            .I(N__33104));
    InMux I__7457 (
            .O(N__33127),
            .I(N__33097));
    InMux I__7456 (
            .O(N__33126),
            .I(N__33094));
    LocalMux I__7455 (
            .O(N__33121),
            .I(N__33091));
    InMux I__7454 (
            .O(N__33120),
            .I(N__33088));
    LocalMux I__7453 (
            .O(N__33117),
            .I(N__33085));
    InMux I__7452 (
            .O(N__33116),
            .I(N__33074));
    InMux I__7451 (
            .O(N__33115),
            .I(N__33074));
    InMux I__7450 (
            .O(N__33114),
            .I(N__33074));
    InMux I__7449 (
            .O(N__33113),
            .I(N__33074));
    InMux I__7448 (
            .O(N__33112),
            .I(N__33074));
    InMux I__7447 (
            .O(N__33111),
            .I(N__33069));
    InMux I__7446 (
            .O(N__33110),
            .I(N__33069));
    InMux I__7445 (
            .O(N__33109),
            .I(N__33066));
    LocalMux I__7444 (
            .O(N__33104),
            .I(N__33063));
    InMux I__7443 (
            .O(N__33103),
            .I(N__33054));
    InMux I__7442 (
            .O(N__33102),
            .I(N__33054));
    InMux I__7441 (
            .O(N__33101),
            .I(N__33054));
    InMux I__7440 (
            .O(N__33100),
            .I(N__33054));
    LocalMux I__7439 (
            .O(N__33097),
            .I(N__33049));
    LocalMux I__7438 (
            .O(N__33094),
            .I(N__33039));
    Span4Mux_v I__7437 (
            .O(N__33091),
            .I(N__33039));
    LocalMux I__7436 (
            .O(N__33088),
            .I(N__33030));
    Span4Mux_h I__7435 (
            .O(N__33085),
            .I(N__33030));
    LocalMux I__7434 (
            .O(N__33074),
            .I(N__33030));
    LocalMux I__7433 (
            .O(N__33069),
            .I(N__33030));
    LocalMux I__7432 (
            .O(N__33066),
            .I(N__33027));
    Span4Mux_v I__7431 (
            .O(N__33063),
            .I(N__33022));
    LocalMux I__7430 (
            .O(N__33054),
            .I(N__33022));
    CascadeMux I__7429 (
            .O(N__33053),
            .I(N__33019));
    CascadeMux I__7428 (
            .O(N__33052),
            .I(N__33016));
    Span4Mux_h I__7427 (
            .O(N__33049),
            .I(N__33009));
    InMux I__7426 (
            .O(N__33048),
            .I(N__33000));
    InMux I__7425 (
            .O(N__33047),
            .I(N__33000));
    InMux I__7424 (
            .O(N__33046),
            .I(N__33000));
    InMux I__7423 (
            .O(N__33045),
            .I(N__33000));
    InMux I__7422 (
            .O(N__33044),
            .I(N__32997));
    Span4Mux_h I__7421 (
            .O(N__33039),
            .I(N__32992));
    Span4Mux_v I__7420 (
            .O(N__33030),
            .I(N__32992));
    Span4Mux_v I__7419 (
            .O(N__33027),
            .I(N__32987));
    Span4Mux_h I__7418 (
            .O(N__33022),
            .I(N__32987));
    InMux I__7417 (
            .O(N__33019),
            .I(N__32974));
    InMux I__7416 (
            .O(N__33016),
            .I(N__32974));
    InMux I__7415 (
            .O(N__33015),
            .I(N__32974));
    InMux I__7414 (
            .O(N__33014),
            .I(N__32974));
    InMux I__7413 (
            .O(N__33013),
            .I(N__32974));
    InMux I__7412 (
            .O(N__33012),
            .I(N__32974));
    Span4Mux_h I__7411 (
            .O(N__33009),
            .I(N__32969));
    LocalMux I__7410 (
            .O(N__33000),
            .I(N__32969));
    LocalMux I__7409 (
            .O(N__32997),
            .I(quadWriteZ0Z_0));
    Odrv4 I__7408 (
            .O(N__32992),
            .I(quadWriteZ0Z_0));
    Odrv4 I__7407 (
            .O(N__32987),
            .I(quadWriteZ0Z_0));
    LocalMux I__7406 (
            .O(N__32974),
            .I(quadWriteZ0Z_0));
    Odrv4 I__7405 (
            .O(N__32969),
            .I(quadWriteZ0Z_0));
    InMux I__7404 (
            .O(N__32958),
            .I(N__32955));
    LocalMux I__7403 (
            .O(N__32955),
            .I(N__32952));
    Odrv12 I__7402 (
            .O(N__32952),
            .I(MOSIrZ0Z_0));
    InMux I__7401 (
            .O(N__32949),
            .I(N__32941));
    InMux I__7400 (
            .O(N__32948),
            .I(N__32938));
    InMux I__7399 (
            .O(N__32947),
            .I(N__32935));
    InMux I__7398 (
            .O(N__32946),
            .I(N__32930));
    InMux I__7397 (
            .O(N__32945),
            .I(N__32930));
    InMux I__7396 (
            .O(N__32944),
            .I(N__32927));
    LocalMux I__7395 (
            .O(N__32941),
            .I(N__32923));
    LocalMux I__7394 (
            .O(N__32938),
            .I(N__32919));
    LocalMux I__7393 (
            .O(N__32935),
            .I(N__32916));
    LocalMux I__7392 (
            .O(N__32930),
            .I(N__32911));
    LocalMux I__7391 (
            .O(N__32927),
            .I(N__32911));
    InMux I__7390 (
            .O(N__32926),
            .I(N__32905));
    Span4Mux_v I__7389 (
            .O(N__32923),
            .I(N__32902));
    InMux I__7388 (
            .O(N__32922),
            .I(N__32899));
    Span4Mux_h I__7387 (
            .O(N__32919),
            .I(N__32892));
    Span4Mux_h I__7386 (
            .O(N__32916),
            .I(N__32892));
    Span4Mux_h I__7385 (
            .O(N__32911),
            .I(N__32892));
    InMux I__7384 (
            .O(N__32910),
            .I(N__32887));
    InMux I__7383 (
            .O(N__32909),
            .I(N__32887));
    InMux I__7382 (
            .O(N__32908),
            .I(N__32884));
    LocalMux I__7381 (
            .O(N__32905),
            .I(data_received_0_repZ0Z2));
    Odrv4 I__7380 (
            .O(N__32902),
            .I(data_received_0_repZ0Z2));
    LocalMux I__7379 (
            .O(N__32899),
            .I(data_received_0_repZ0Z2));
    Odrv4 I__7378 (
            .O(N__32892),
            .I(data_received_0_repZ0Z2));
    LocalMux I__7377 (
            .O(N__32887),
            .I(data_received_0_repZ0Z2));
    LocalMux I__7376 (
            .O(N__32884),
            .I(data_received_0_repZ0Z2));
    InMux I__7375 (
            .O(N__32871),
            .I(N__32868));
    LocalMux I__7374 (
            .O(N__32868),
            .I(N__32863));
    InMux I__7373 (
            .O(N__32867),
            .I(N__32860));
    InMux I__7372 (
            .O(N__32866),
            .I(N__32857));
    Span4Mux_v I__7371 (
            .O(N__32863),
            .I(N__32854));
    LocalMux I__7370 (
            .O(N__32860),
            .I(N__32851));
    LocalMux I__7369 (
            .O(N__32857),
            .I(N__32848));
    Odrv4 I__7368 (
            .O(N__32854),
            .I(dataRead4_10));
    Odrv4 I__7367 (
            .O(N__32851),
            .I(dataRead4_10));
    Odrv4 I__7366 (
            .O(N__32848),
            .I(dataRead4_10));
    CascadeMux I__7365 (
            .O(N__32841),
            .I(N__32836));
    CascadeMux I__7364 (
            .O(N__32840),
            .I(N__32832));
    InMux I__7363 (
            .O(N__32839),
            .I(N__32827));
    InMux I__7362 (
            .O(N__32836),
            .I(N__32822));
    InMux I__7361 (
            .O(N__32835),
            .I(N__32822));
    InMux I__7360 (
            .O(N__32832),
            .I(N__32819));
    InMux I__7359 (
            .O(N__32831),
            .I(N__32815));
    InMux I__7358 (
            .O(N__32830),
            .I(N__32812));
    LocalMux I__7357 (
            .O(N__32827),
            .I(N__32807));
    LocalMux I__7356 (
            .O(N__32822),
            .I(N__32802));
    LocalMux I__7355 (
            .O(N__32819),
            .I(N__32802));
    CascadeMux I__7354 (
            .O(N__32818),
            .I(N__32797));
    LocalMux I__7353 (
            .O(N__32815),
            .I(N__32794));
    LocalMux I__7352 (
            .O(N__32812),
            .I(N__32791));
    InMux I__7351 (
            .O(N__32811),
            .I(N__32788));
    InMux I__7350 (
            .O(N__32810),
            .I(N__32785));
    Span4Mux_h I__7349 (
            .O(N__32807),
            .I(N__32780));
    Span4Mux_h I__7348 (
            .O(N__32802),
            .I(N__32780));
    InMux I__7347 (
            .O(N__32801),
            .I(N__32775));
    InMux I__7346 (
            .O(N__32800),
            .I(N__32775));
    InMux I__7345 (
            .O(N__32797),
            .I(N__32772));
    Odrv4 I__7344 (
            .O(N__32794),
            .I(data_received_2_repZ0Z2));
    Odrv4 I__7343 (
            .O(N__32791),
            .I(data_received_2_repZ0Z2));
    LocalMux I__7342 (
            .O(N__32788),
            .I(data_received_2_repZ0Z2));
    LocalMux I__7341 (
            .O(N__32785),
            .I(data_received_2_repZ0Z2));
    Odrv4 I__7340 (
            .O(N__32780),
            .I(data_received_2_repZ0Z2));
    LocalMux I__7339 (
            .O(N__32775),
            .I(data_received_2_repZ0Z2));
    LocalMux I__7338 (
            .O(N__32772),
            .I(data_received_2_repZ0Z2));
    InMux I__7337 (
            .O(N__32757),
            .I(N__32754));
    LocalMux I__7336 (
            .O(N__32754),
            .I(\QuadInstance0.Quad_RNO_0_0_10 ));
    InMux I__7335 (
            .O(N__32751),
            .I(N__32747));
    InMux I__7334 (
            .O(N__32750),
            .I(N__32744));
    LocalMux I__7333 (
            .O(N__32747),
            .I(\QuadInstance0.delayedCh_BZ0Z_1 ));
    LocalMux I__7332 (
            .O(N__32744),
            .I(\QuadInstance0.delayedCh_BZ0Z_1 ));
    InMux I__7331 (
            .O(N__32739),
            .I(N__32736));
    LocalMux I__7330 (
            .O(N__32736),
            .I(\QuadInstance0.delayedCh_AZ0Z_2 ));
    InMux I__7329 (
            .O(N__32733),
            .I(N__32730));
    LocalMux I__7328 (
            .O(N__32730),
            .I(N__32726));
    InMux I__7327 (
            .O(N__32729),
            .I(N__32723));
    Span4Mux_v I__7326 (
            .O(N__32726),
            .I(N__32720));
    LocalMux I__7325 (
            .O(N__32723),
            .I(N__32717));
    Span4Mux_h I__7324 (
            .O(N__32720),
            .I(N__32713));
    Span4Mux_v I__7323 (
            .O(N__32717),
            .I(N__32710));
    InMux I__7322 (
            .O(N__32716),
            .I(N__32707));
    Odrv4 I__7321 (
            .O(N__32713),
            .I(dataRead0_1));
    Odrv4 I__7320 (
            .O(N__32710),
            .I(dataRead0_1));
    LocalMux I__7319 (
            .O(N__32707),
            .I(dataRead0_1));
    CascadeMux I__7318 (
            .O(N__32700),
            .I(\QuadInstance0.count_enable_cascade_ ));
    CascadeMux I__7317 (
            .O(N__32697),
            .I(N__32694));
    InMux I__7316 (
            .O(N__32694),
            .I(N__32691));
    LocalMux I__7315 (
            .O(N__32691),
            .I(\QuadInstance0.Quad_RNIGEBH1Z0Z_1 ));
    CascadeMux I__7314 (
            .O(N__32688),
            .I(N__32684));
    InMux I__7313 (
            .O(N__32687),
            .I(N__32680));
    InMux I__7312 (
            .O(N__32684),
            .I(N__32675));
    InMux I__7311 (
            .O(N__32683),
            .I(N__32675));
    LocalMux I__7310 (
            .O(N__32680),
            .I(dataRead0_10));
    LocalMux I__7309 (
            .O(N__32675),
            .I(dataRead0_10));
    CascadeMux I__7308 (
            .O(N__32670),
            .I(N__32667));
    InMux I__7307 (
            .O(N__32667),
            .I(N__32664));
    LocalMux I__7306 (
            .O(N__32664),
            .I(\QuadInstance0.Quad_RNI0L8Q1Z0Z_10 ));
    InMux I__7305 (
            .O(N__32661),
            .I(N__32658));
    LocalMux I__7304 (
            .O(N__32658),
            .I(N__32654));
    InMux I__7303 (
            .O(N__32657),
            .I(N__32651));
    Span4Mux_h I__7302 (
            .O(N__32654),
            .I(N__32645));
    LocalMux I__7301 (
            .O(N__32651),
            .I(N__32645));
    InMux I__7300 (
            .O(N__32650),
            .I(N__32642));
    Odrv4 I__7299 (
            .O(N__32645),
            .I(dataRead0_2));
    LocalMux I__7298 (
            .O(N__32642),
            .I(dataRead0_2));
    CascadeMux I__7297 (
            .O(N__32637),
            .I(N__32634));
    InMux I__7296 (
            .O(N__32634),
            .I(N__32631));
    LocalMux I__7295 (
            .O(N__32631),
            .I(\QuadInstance0.Quad_RNIHFBH1Z0Z_2 ));
    InMux I__7294 (
            .O(N__32628),
            .I(N__32622));
    InMux I__7293 (
            .O(N__32627),
            .I(N__32622));
    LocalMux I__7292 (
            .O(N__32622),
            .I(\QuadInstance0.delayedCh_BZ0Z_2 ));
    CascadeMux I__7291 (
            .O(N__32619),
            .I(N__32616));
    InMux I__7290 (
            .O(N__32616),
            .I(N__32613));
    LocalMux I__7289 (
            .O(N__32613),
            .I(N__32610));
    Odrv4 I__7288 (
            .O(N__32610),
            .I(\PWMInstance2.un1_PWMPulseWidthCount_0_I_27_c_RNO_1 ));
    InMux I__7287 (
            .O(N__32607),
            .I(N__32604));
    LocalMux I__7286 (
            .O(N__32604),
            .I(N__32601));
    Odrv4 I__7285 (
            .O(N__32601),
            .I(\PWMInstance2.un1_PWMPulseWidthCount_0_I_45_c_RNO_1 ));
    InMux I__7284 (
            .O(N__32598),
            .I(N__32595));
    LocalMux I__7283 (
            .O(N__32595),
            .I(\PWMInstance2.un1_PWMPulseWidthCount_0_I_39_c_RNO_1 ));
    CascadeMux I__7282 (
            .O(N__32592),
            .I(N__32563));
    CascadeMux I__7281 (
            .O(N__32591),
            .I(N__32560));
    CascadeMux I__7280 (
            .O(N__32590),
            .I(N__32557));
    CascadeMux I__7279 (
            .O(N__32589),
            .I(N__32554));
    CascadeMux I__7278 (
            .O(N__32588),
            .I(N__32551));
    CascadeMux I__7277 (
            .O(N__32587),
            .I(N__32548));
    CascadeMux I__7276 (
            .O(N__32586),
            .I(N__32545));
    CascadeMux I__7275 (
            .O(N__32585),
            .I(N__32535));
    CascadeMux I__7274 (
            .O(N__32584),
            .I(N__32531));
    CascadeMux I__7273 (
            .O(N__32583),
            .I(N__32528));
    CascadeMux I__7272 (
            .O(N__32582),
            .I(N__32525));
    CascadeMux I__7271 (
            .O(N__32581),
            .I(N__32522));
    CascadeMux I__7270 (
            .O(N__32580),
            .I(N__32519));
    CascadeMux I__7269 (
            .O(N__32579),
            .I(N__32515));
    CascadeMux I__7268 (
            .O(N__32578),
            .I(N__32512));
    CascadeMux I__7267 (
            .O(N__32577),
            .I(N__32509));
    CascadeMux I__7266 (
            .O(N__32576),
            .I(N__32506));
    CascadeMux I__7265 (
            .O(N__32575),
            .I(N__32503));
    CascadeMux I__7264 (
            .O(N__32574),
            .I(N__32500));
    CascadeMux I__7263 (
            .O(N__32573),
            .I(N__32497));
    CascadeMux I__7262 (
            .O(N__32572),
            .I(N__32491));
    CascadeMux I__7261 (
            .O(N__32571),
            .I(N__32488));
    CascadeMux I__7260 (
            .O(N__32570),
            .I(N__32485));
    CascadeMux I__7259 (
            .O(N__32569),
            .I(N__32482));
    CascadeMux I__7258 (
            .O(N__32568),
            .I(N__32479));
    CascadeMux I__7257 (
            .O(N__32567),
            .I(N__32476));
    CascadeMux I__7256 (
            .O(N__32566),
            .I(N__32473));
    InMux I__7255 (
            .O(N__32563),
            .I(N__32457));
    InMux I__7254 (
            .O(N__32560),
            .I(N__32457));
    InMux I__7253 (
            .O(N__32557),
            .I(N__32457));
    InMux I__7252 (
            .O(N__32554),
            .I(N__32457));
    InMux I__7251 (
            .O(N__32551),
            .I(N__32450));
    InMux I__7250 (
            .O(N__32548),
            .I(N__32450));
    InMux I__7249 (
            .O(N__32545),
            .I(N__32450));
    CascadeMux I__7248 (
            .O(N__32544),
            .I(N__32447));
    CascadeMux I__7247 (
            .O(N__32543),
            .I(N__32444));
    CascadeMux I__7246 (
            .O(N__32542),
            .I(N__32441));
    CascadeMux I__7245 (
            .O(N__32541),
            .I(N__32438));
    CascadeMux I__7244 (
            .O(N__32540),
            .I(N__32435));
    CascadeMux I__7243 (
            .O(N__32539),
            .I(N__32432));
    CascadeMux I__7242 (
            .O(N__32538),
            .I(N__32429));
    InMux I__7241 (
            .O(N__32535),
            .I(N__32418));
    InMux I__7240 (
            .O(N__32534),
            .I(N__32418));
    InMux I__7239 (
            .O(N__32531),
            .I(N__32418));
    InMux I__7238 (
            .O(N__32528),
            .I(N__32418));
    InMux I__7237 (
            .O(N__32525),
            .I(N__32418));
    InMux I__7236 (
            .O(N__32522),
            .I(N__32413));
    InMux I__7235 (
            .O(N__32519),
            .I(N__32413));
    CascadeMux I__7234 (
            .O(N__32518),
            .I(N__32407));
    InMux I__7233 (
            .O(N__32515),
            .I(N__32398));
    InMux I__7232 (
            .O(N__32512),
            .I(N__32398));
    InMux I__7231 (
            .O(N__32509),
            .I(N__32398));
    InMux I__7230 (
            .O(N__32506),
            .I(N__32398));
    InMux I__7229 (
            .O(N__32503),
            .I(N__32391));
    InMux I__7228 (
            .O(N__32500),
            .I(N__32391));
    InMux I__7227 (
            .O(N__32497),
            .I(N__32391));
    CascadeMux I__7226 (
            .O(N__32496),
            .I(N__32387));
    CascadeMux I__7225 (
            .O(N__32495),
            .I(N__32384));
    CascadeMux I__7224 (
            .O(N__32494),
            .I(N__32379));
    InMux I__7223 (
            .O(N__32491),
            .I(N__32370));
    InMux I__7222 (
            .O(N__32488),
            .I(N__32370));
    InMux I__7221 (
            .O(N__32485),
            .I(N__32370));
    InMux I__7220 (
            .O(N__32482),
            .I(N__32370));
    InMux I__7219 (
            .O(N__32479),
            .I(N__32363));
    InMux I__7218 (
            .O(N__32476),
            .I(N__32363));
    InMux I__7217 (
            .O(N__32473),
            .I(N__32363));
    CascadeMux I__7216 (
            .O(N__32472),
            .I(N__32360));
    CascadeMux I__7215 (
            .O(N__32471),
            .I(N__32357));
    CascadeMux I__7214 (
            .O(N__32470),
            .I(N__32354));
    CascadeMux I__7213 (
            .O(N__32469),
            .I(N__32351));
    CascadeMux I__7212 (
            .O(N__32468),
            .I(N__32348));
    CascadeMux I__7211 (
            .O(N__32467),
            .I(N__32345));
    CascadeMux I__7210 (
            .O(N__32466),
            .I(N__32342));
    LocalMux I__7209 (
            .O(N__32457),
            .I(N__32339));
    LocalMux I__7208 (
            .O(N__32450),
            .I(N__32336));
    InMux I__7207 (
            .O(N__32447),
            .I(N__32327));
    InMux I__7206 (
            .O(N__32444),
            .I(N__32327));
    InMux I__7205 (
            .O(N__32441),
            .I(N__32327));
    InMux I__7204 (
            .O(N__32438),
            .I(N__32327));
    InMux I__7203 (
            .O(N__32435),
            .I(N__32320));
    InMux I__7202 (
            .O(N__32432),
            .I(N__32320));
    InMux I__7201 (
            .O(N__32429),
            .I(N__32320));
    LocalMux I__7200 (
            .O(N__32418),
            .I(N__32315));
    LocalMux I__7199 (
            .O(N__32413),
            .I(N__32315));
    CascadeMux I__7198 (
            .O(N__32412),
            .I(N__32311));
    CascadeMux I__7197 (
            .O(N__32411),
            .I(N__32308));
    CascadeMux I__7196 (
            .O(N__32410),
            .I(N__32302));
    InMux I__7195 (
            .O(N__32407),
            .I(N__32299));
    LocalMux I__7194 (
            .O(N__32398),
            .I(N__32294));
    LocalMux I__7193 (
            .O(N__32391),
            .I(N__32294));
    InMux I__7192 (
            .O(N__32390),
            .I(N__32281));
    InMux I__7191 (
            .O(N__32387),
            .I(N__32281));
    InMux I__7190 (
            .O(N__32384),
            .I(N__32281));
    InMux I__7189 (
            .O(N__32383),
            .I(N__32281));
    InMux I__7188 (
            .O(N__32382),
            .I(N__32281));
    InMux I__7187 (
            .O(N__32379),
            .I(N__32281));
    LocalMux I__7186 (
            .O(N__32370),
            .I(N__32276));
    LocalMux I__7185 (
            .O(N__32363),
            .I(N__32276));
    InMux I__7184 (
            .O(N__32360),
            .I(N__32267));
    InMux I__7183 (
            .O(N__32357),
            .I(N__32267));
    InMux I__7182 (
            .O(N__32354),
            .I(N__32267));
    InMux I__7181 (
            .O(N__32351),
            .I(N__32267));
    InMux I__7180 (
            .O(N__32348),
            .I(N__32260));
    InMux I__7179 (
            .O(N__32345),
            .I(N__32260));
    InMux I__7178 (
            .O(N__32342),
            .I(N__32260));
    Span4Mux_v I__7177 (
            .O(N__32339),
            .I(N__32255));
    Span4Mux_v I__7176 (
            .O(N__32336),
            .I(N__32255));
    LocalMux I__7175 (
            .O(N__32327),
            .I(N__32250));
    LocalMux I__7174 (
            .O(N__32320),
            .I(N__32250));
    Span4Mux_v I__7173 (
            .O(N__32315),
            .I(N__32247));
    InMux I__7172 (
            .O(N__32314),
            .I(N__32232));
    InMux I__7171 (
            .O(N__32311),
            .I(N__32232));
    InMux I__7170 (
            .O(N__32308),
            .I(N__32232));
    InMux I__7169 (
            .O(N__32307),
            .I(N__32232));
    InMux I__7168 (
            .O(N__32306),
            .I(N__32232));
    InMux I__7167 (
            .O(N__32305),
            .I(N__32232));
    InMux I__7166 (
            .O(N__32302),
            .I(N__32232));
    LocalMux I__7165 (
            .O(N__32299),
            .I(N__32229));
    Span4Mux_h I__7164 (
            .O(N__32294),
            .I(N__32224));
    LocalMux I__7163 (
            .O(N__32281),
            .I(N__32224));
    Span4Mux_h I__7162 (
            .O(N__32276),
            .I(N__32221));
    LocalMux I__7161 (
            .O(N__32267),
            .I(N__32216));
    LocalMux I__7160 (
            .O(N__32260),
            .I(N__32216));
    Span4Mux_h I__7159 (
            .O(N__32255),
            .I(N__32211));
    Span4Mux_h I__7158 (
            .O(N__32250),
            .I(N__32211));
    Sp12to4 I__7157 (
            .O(N__32247),
            .I(N__32208));
    LocalMux I__7156 (
            .O(N__32232),
            .I(N__32205));
    Span4Mux_v I__7155 (
            .O(N__32229),
            .I(N__32202));
    Span4Mux_v I__7154 (
            .O(N__32224),
            .I(N__32199));
    Span4Mux_v I__7153 (
            .O(N__32221),
            .I(N__32194));
    Span4Mux_h I__7152 (
            .O(N__32216),
            .I(N__32194));
    Span4Mux_v I__7151 (
            .O(N__32211),
            .I(N__32191));
    Span12Mux_h I__7150 (
            .O(N__32208),
            .I(N__32186));
    Sp12to4 I__7149 (
            .O(N__32205),
            .I(N__32186));
    Span4Mux_h I__7148 (
            .O(N__32202),
            .I(N__32179));
    Span4Mux_h I__7147 (
            .O(N__32199),
            .I(N__32179));
    Span4Mux_h I__7146 (
            .O(N__32194),
            .I(N__32179));
    Odrv4 I__7145 (
            .O(N__32191),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__7144 (
            .O(N__32186),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__7143 (
            .O(N__32179),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__7142 (
            .O(N__32172),
            .I(N__32169));
    InMux I__7141 (
            .O(N__32169),
            .I(N__32166));
    LocalMux I__7140 (
            .O(N__32166),
            .I(\PWMInstance2.un1_PWMPulseWidthCount_0_I_21_c_RNO_1 ));
    InMux I__7139 (
            .O(N__32163),
            .I(N__32160));
    LocalMux I__7138 (
            .O(N__32160),
            .I(N__32157));
    Odrv12 I__7137 (
            .O(N__32157),
            .I(\PWMInstance2.un1_periodCounter12_1_0_a2_0 ));
    InMux I__7136 (
            .O(N__32154),
            .I(bfn_17_15_0_));
    IoInMux I__7135 (
            .O(N__32151),
            .I(N__32148));
    LocalMux I__7134 (
            .O(N__32148),
            .I(N__32145));
    Span4Mux_s1_v I__7133 (
            .O(N__32145),
            .I(N__32142));
    Span4Mux_v I__7132 (
            .O(N__32142),
            .I(N__32138));
    InMux I__7131 (
            .O(N__32141),
            .I(N__32135));
    Odrv4 I__7130 (
            .O(N__32138),
            .I(PWM2_c));
    LocalMux I__7129 (
            .O(N__32135),
            .I(PWM2_c));
    InMux I__7128 (
            .O(N__32130),
            .I(N__32127));
    LocalMux I__7127 (
            .O(N__32127),
            .I(MOSI_c));
    InMux I__7126 (
            .O(N__32124),
            .I(N__32121));
    LocalMux I__7125 (
            .O(N__32121),
            .I(ch1_A_c));
    InMux I__7124 (
            .O(N__32118),
            .I(N__32115));
    LocalMux I__7123 (
            .O(N__32115),
            .I(N__32112));
    Span4Mux_h I__7122 (
            .O(N__32112),
            .I(N__32109));
    Odrv4 I__7121 (
            .O(N__32109),
            .I(\QuadInstance1.delayedCh_AZ0Z_0 ));
    InMux I__7120 (
            .O(N__32106),
            .I(N__32103));
    LocalMux I__7119 (
            .O(N__32103),
            .I(N__32100));
    Span4Mux_h I__7118 (
            .O(N__32100),
            .I(N__32097));
    Span4Mux_h I__7117 (
            .O(N__32097),
            .I(N__32094));
    Odrv4 I__7116 (
            .O(N__32094),
            .I(\QuadInstance0.delayedCh_AZ0Z_0 ));
    InMux I__7115 (
            .O(N__32091),
            .I(N__32088));
    LocalMux I__7114 (
            .O(N__32088),
            .I(N__32079));
    InMux I__7113 (
            .O(N__32087),
            .I(N__32074));
    InMux I__7112 (
            .O(N__32086),
            .I(N__32074));
    InMux I__7111 (
            .O(N__32085),
            .I(N__32069));
    InMux I__7110 (
            .O(N__32084),
            .I(N__32066));
    InMux I__7109 (
            .O(N__32083),
            .I(N__32063));
    InMux I__7108 (
            .O(N__32082),
            .I(N__32060));
    Span4Mux_v I__7107 (
            .O(N__32079),
            .I(N__32057));
    LocalMux I__7106 (
            .O(N__32074),
            .I(N__32054));
    InMux I__7105 (
            .O(N__32073),
            .I(N__32051));
    InMux I__7104 (
            .O(N__32072),
            .I(N__32047));
    LocalMux I__7103 (
            .O(N__32069),
            .I(N__32044));
    LocalMux I__7102 (
            .O(N__32066),
            .I(N__32040));
    LocalMux I__7101 (
            .O(N__32063),
            .I(N__32037));
    LocalMux I__7100 (
            .O(N__32060),
            .I(N__32034));
    Span4Mux_h I__7099 (
            .O(N__32057),
            .I(N__32026));
    Span4Mux_v I__7098 (
            .O(N__32054),
            .I(N__32026));
    LocalMux I__7097 (
            .O(N__32051),
            .I(N__32026));
    InMux I__7096 (
            .O(N__32050),
            .I(N__32023));
    LocalMux I__7095 (
            .O(N__32047),
            .I(N__32017));
    Span4Mux_h I__7094 (
            .O(N__32044),
            .I(N__32014));
    InMux I__7093 (
            .O(N__32043),
            .I(N__32011));
    Span4Mux_h I__7092 (
            .O(N__32040),
            .I(N__32008));
    Span4Mux_h I__7091 (
            .O(N__32037),
            .I(N__32005));
    Span4Mux_v I__7090 (
            .O(N__32034),
            .I(N__32002));
    InMux I__7089 (
            .O(N__32033),
            .I(N__31999));
    Span4Mux_h I__7088 (
            .O(N__32026),
            .I(N__31994));
    LocalMux I__7087 (
            .O(N__32023),
            .I(N__31994));
    InMux I__7086 (
            .O(N__32022),
            .I(N__31989));
    InMux I__7085 (
            .O(N__32021),
            .I(N__31989));
    InMux I__7084 (
            .O(N__32020),
            .I(N__31986));
    Span4Mux_h I__7083 (
            .O(N__32017),
            .I(N__31978));
    Span4Mux_h I__7082 (
            .O(N__32014),
            .I(N__31978));
    LocalMux I__7081 (
            .O(N__32011),
            .I(N__31978));
    Span4Mux_h I__7080 (
            .O(N__32008),
            .I(N__31973));
    Span4Mux_v I__7079 (
            .O(N__32005),
            .I(N__31973));
    Span4Mux_h I__7078 (
            .O(N__32002),
            .I(N__31970));
    LocalMux I__7077 (
            .O(N__31999),
            .I(N__31967));
    Span4Mux_v I__7076 (
            .O(N__31994),
            .I(N__31964));
    LocalMux I__7075 (
            .O(N__31989),
            .I(N__31959));
    LocalMux I__7074 (
            .O(N__31986),
            .I(N__31959));
    InMux I__7073 (
            .O(N__31985),
            .I(N__31956));
    Span4Mux_v I__7072 (
            .O(N__31978),
            .I(N__31951));
    Span4Mux_h I__7071 (
            .O(N__31973),
            .I(N__31951));
    Span4Mux_h I__7070 (
            .O(N__31970),
            .I(N__31942));
    Span4Mux_h I__7069 (
            .O(N__31967),
            .I(N__31942));
    Span4Mux_h I__7068 (
            .O(N__31964),
            .I(N__31942));
    Span4Mux_h I__7067 (
            .O(N__31959),
            .I(N__31942));
    LocalMux I__7066 (
            .O(N__31956),
            .I(dataWriteZ0Z_3));
    Odrv4 I__7065 (
            .O(N__31951),
            .I(dataWriteZ0Z_3));
    Odrv4 I__7064 (
            .O(N__31942),
            .I(dataWriteZ0Z_3));
    InMux I__7063 (
            .O(N__31935),
            .I(N__31932));
    LocalMux I__7062 (
            .O(N__31932),
            .I(\PWMInstance2.PWMPulseWidthCountZ0Z_3 ));
    InMux I__7061 (
            .O(N__31929),
            .I(N__31926));
    LocalMux I__7060 (
            .O(N__31926),
            .I(\PWMInstance2.PWMPulseWidthCountZ0Z_14 ));
    CascadeMux I__7059 (
            .O(N__31923),
            .I(N__31920));
    InMux I__7058 (
            .O(N__31920),
            .I(N__31913));
    CascadeMux I__7057 (
            .O(N__31919),
            .I(N__31910));
    InMux I__7056 (
            .O(N__31918),
            .I(N__31905));
    CascadeMux I__7055 (
            .O(N__31917),
            .I(N__31900));
    CascadeMux I__7054 (
            .O(N__31916),
            .I(N__31897));
    LocalMux I__7053 (
            .O(N__31913),
            .I(N__31891));
    InMux I__7052 (
            .O(N__31910),
            .I(N__31888));
    CascadeMux I__7051 (
            .O(N__31909),
            .I(N__31885));
    CascadeMux I__7050 (
            .O(N__31908),
            .I(N__31882));
    LocalMux I__7049 (
            .O(N__31905),
            .I(N__31879));
    InMux I__7048 (
            .O(N__31904),
            .I(N__31875));
    InMux I__7047 (
            .O(N__31903),
            .I(N__31872));
    InMux I__7046 (
            .O(N__31900),
            .I(N__31868));
    InMux I__7045 (
            .O(N__31897),
            .I(N__31865));
    CascadeMux I__7044 (
            .O(N__31896),
            .I(N__31862));
    CascadeMux I__7043 (
            .O(N__31895),
            .I(N__31859));
    InMux I__7042 (
            .O(N__31894),
            .I(N__31854));
    Span4Mux_h I__7041 (
            .O(N__31891),
            .I(N__31849));
    LocalMux I__7040 (
            .O(N__31888),
            .I(N__31849));
    InMux I__7039 (
            .O(N__31885),
            .I(N__31846));
    InMux I__7038 (
            .O(N__31882),
            .I(N__31843));
    Span4Mux_v I__7037 (
            .O(N__31879),
            .I(N__31840));
    InMux I__7036 (
            .O(N__31878),
            .I(N__31837));
    LocalMux I__7035 (
            .O(N__31875),
            .I(N__31832));
    LocalMux I__7034 (
            .O(N__31872),
            .I(N__31832));
    InMux I__7033 (
            .O(N__31871),
            .I(N__31829));
    LocalMux I__7032 (
            .O(N__31868),
            .I(N__31826));
    LocalMux I__7031 (
            .O(N__31865),
            .I(N__31823));
    InMux I__7030 (
            .O(N__31862),
            .I(N__31820));
    InMux I__7029 (
            .O(N__31859),
            .I(N__31817));
    InMux I__7028 (
            .O(N__31858),
            .I(N__31814));
    InMux I__7027 (
            .O(N__31857),
            .I(N__31811));
    LocalMux I__7026 (
            .O(N__31854),
            .I(N__31808));
    Span4Mux_v I__7025 (
            .O(N__31849),
            .I(N__31801));
    LocalMux I__7024 (
            .O(N__31846),
            .I(N__31801));
    LocalMux I__7023 (
            .O(N__31843),
            .I(N__31801));
    Span4Mux_h I__7022 (
            .O(N__31840),
            .I(N__31798));
    LocalMux I__7021 (
            .O(N__31837),
            .I(N__31795));
    Span4Mux_v I__7020 (
            .O(N__31832),
            .I(N__31792));
    LocalMux I__7019 (
            .O(N__31829),
            .I(N__31789));
    Span4Mux_v I__7018 (
            .O(N__31826),
            .I(N__31786));
    Span4Mux_h I__7017 (
            .O(N__31823),
            .I(N__31779));
    LocalMux I__7016 (
            .O(N__31820),
            .I(N__31779));
    LocalMux I__7015 (
            .O(N__31817),
            .I(N__31779));
    LocalMux I__7014 (
            .O(N__31814),
            .I(N__31776));
    LocalMux I__7013 (
            .O(N__31811),
            .I(N__31773));
    Span4Mux_v I__7012 (
            .O(N__31808),
            .I(N__31768));
    Span4Mux_v I__7011 (
            .O(N__31801),
            .I(N__31768));
    Span4Mux_v I__7010 (
            .O(N__31798),
            .I(N__31765));
    Span4Mux_v I__7009 (
            .O(N__31795),
            .I(N__31758));
    Span4Mux_h I__7008 (
            .O(N__31792),
            .I(N__31758));
    Span4Mux_v I__7007 (
            .O(N__31789),
            .I(N__31758));
    Span4Mux_h I__7006 (
            .O(N__31786),
            .I(N__31753));
    Span4Mux_v I__7005 (
            .O(N__31779),
            .I(N__31753));
    Span4Mux_v I__7004 (
            .O(N__31776),
            .I(N__31746));
    Span4Mux_v I__7003 (
            .O(N__31773),
            .I(N__31746));
    Span4Mux_h I__7002 (
            .O(N__31768),
            .I(N__31746));
    Odrv4 I__7001 (
            .O(N__31765),
            .I(dataWriteZ0Z_15));
    Odrv4 I__7000 (
            .O(N__31758),
            .I(dataWriteZ0Z_15));
    Odrv4 I__6999 (
            .O(N__31753),
            .I(dataWriteZ0Z_15));
    Odrv4 I__6998 (
            .O(N__31746),
            .I(dataWriteZ0Z_15));
    InMux I__6997 (
            .O(N__31737),
            .I(N__31734));
    LocalMux I__6996 (
            .O(N__31734),
            .I(\PWMInstance2.PWMPulseWidthCountZ0Z_15 ));
    InMux I__6995 (
            .O(N__31731),
            .I(N__31728));
    LocalMux I__6994 (
            .O(N__31728),
            .I(N__31725));
    Span4Mux_h I__6993 (
            .O(N__31725),
            .I(N__31722));
    Odrv4 I__6992 (
            .O(N__31722),
            .I(\PWMInstance2.PWMPulseWidthCountZ0Z_13 ));
    InMux I__6991 (
            .O(N__31719),
            .I(N__31716));
    LocalMux I__6990 (
            .O(N__31716),
            .I(N__31713));
    Odrv4 I__6989 (
            .O(N__31713),
            .I(\PWMInstance2.PWMPulseWidthCountZ0Z_12 ));
    InMux I__6988 (
            .O(N__31710),
            .I(N__31707));
    LocalMux I__6987 (
            .O(N__31707),
            .I(N__31704));
    Odrv12 I__6986 (
            .O(N__31704),
            .I(\PWMInstance2.un1_PWMPulseWidthCount_0_I_1_c_RNO_1 ));
    CascadeMux I__6985 (
            .O(N__31701),
            .I(N__31698));
    InMux I__6984 (
            .O(N__31698),
            .I(N__31695));
    LocalMux I__6983 (
            .O(N__31695),
            .I(\PWMInstance2.un1_PWMPulseWidthCount_0_I_9_c_RNO_1 ));
    InMux I__6982 (
            .O(N__31692),
            .I(N__31683));
    InMux I__6981 (
            .O(N__31691),
            .I(N__31683));
    InMux I__6980 (
            .O(N__31690),
            .I(N__31683));
    LocalMux I__6979 (
            .O(N__31683),
            .I(N__31680));
    Odrv4 I__6978 (
            .O(N__31680),
            .I(pwmWriteZ0Z_2));
    InMux I__6977 (
            .O(N__31677),
            .I(N__31671));
    InMux I__6976 (
            .O(N__31676),
            .I(N__31671));
    LocalMux I__6975 (
            .O(N__31671),
            .I(N__31668));
    Odrv12 I__6974 (
            .O(N__31668),
            .I(pwmWrite_fastZ0Z_2));
    CascadeMux I__6973 (
            .O(N__31665),
            .I(N__31661));
    CascadeMux I__6972 (
            .O(N__31664),
            .I(N__31658));
    InMux I__6971 (
            .O(N__31661),
            .I(N__31647));
    InMux I__6970 (
            .O(N__31658),
            .I(N__31647));
    InMux I__6969 (
            .O(N__31657),
            .I(N__31647));
    InMux I__6968 (
            .O(N__31656),
            .I(N__31647));
    LocalMux I__6967 (
            .O(N__31647),
            .I(\PWMInstance2.clkCountZ0Z_1 ));
    InMux I__6966 (
            .O(N__31644),
            .I(N__31632));
    InMux I__6965 (
            .O(N__31643),
            .I(N__31632));
    InMux I__6964 (
            .O(N__31642),
            .I(N__31632));
    InMux I__6963 (
            .O(N__31641),
            .I(N__31632));
    LocalMux I__6962 (
            .O(N__31632),
            .I(\PWMInstance2.clkCountZ0Z_0 ));
    CascadeMux I__6961 (
            .O(N__31629),
            .I(\PWMInstance2.un1_periodCounter12_1_0_a2_0_6_cascade_ ));
    InMux I__6960 (
            .O(N__31626),
            .I(N__31623));
    LocalMux I__6959 (
            .O(N__31623),
            .I(\PWMInstance2.un1_periodCounter12_1_0_a2_0_9 ));
    CascadeMux I__6958 (
            .O(N__31620),
            .I(\PWMInstance2.un1_periodCounter12_1_0_a2_0_14_cascade_ ));
    InMux I__6957 (
            .O(N__31617),
            .I(N__31614));
    LocalMux I__6956 (
            .O(N__31614),
            .I(N__31611));
    Odrv4 I__6955 (
            .O(N__31611),
            .I(\PWMInstance2.un1_periodCounter12_1_0_a2_0_10 ));
    InMux I__6954 (
            .O(N__31608),
            .I(N__31605));
    LocalMux I__6953 (
            .O(N__31605),
            .I(N__31600));
    InMux I__6952 (
            .O(N__31604),
            .I(N__31597));
    InMux I__6951 (
            .O(N__31603),
            .I(N__31594));
    Span4Mux_s2_v I__6950 (
            .O(N__31600),
            .I(N__31580));
    LocalMux I__6949 (
            .O(N__31597),
            .I(N__31577));
    LocalMux I__6948 (
            .O(N__31594),
            .I(N__31574));
    InMux I__6947 (
            .O(N__31593),
            .I(N__31571));
    InMux I__6946 (
            .O(N__31592),
            .I(N__31568));
    InMux I__6945 (
            .O(N__31591),
            .I(N__31565));
    InMux I__6944 (
            .O(N__31590),
            .I(N__31560));
    InMux I__6943 (
            .O(N__31589),
            .I(N__31560));
    InMux I__6942 (
            .O(N__31588),
            .I(N__31555));
    InMux I__6941 (
            .O(N__31587),
            .I(N__31555));
    InMux I__6940 (
            .O(N__31586),
            .I(N__31550));
    InMux I__6939 (
            .O(N__31585),
            .I(N__31550));
    InMux I__6938 (
            .O(N__31584),
            .I(N__31547));
    InMux I__6937 (
            .O(N__31583),
            .I(N__31544));
    Span4Mux_v I__6936 (
            .O(N__31580),
            .I(N__31539));
    Span4Mux_v I__6935 (
            .O(N__31577),
            .I(N__31534));
    Span4Mux_v I__6934 (
            .O(N__31574),
            .I(N__31534));
    LocalMux I__6933 (
            .O(N__31571),
            .I(N__31531));
    LocalMux I__6932 (
            .O(N__31568),
            .I(N__31528));
    LocalMux I__6931 (
            .O(N__31565),
            .I(N__31525));
    LocalMux I__6930 (
            .O(N__31560),
            .I(N__31520));
    LocalMux I__6929 (
            .O(N__31555),
            .I(N__31520));
    LocalMux I__6928 (
            .O(N__31550),
            .I(N__31517));
    LocalMux I__6927 (
            .O(N__31547),
            .I(N__31512));
    LocalMux I__6926 (
            .O(N__31544),
            .I(N__31512));
    InMux I__6925 (
            .O(N__31543),
            .I(N__31509));
    InMux I__6924 (
            .O(N__31542),
            .I(N__31506));
    Span4Mux_v I__6923 (
            .O(N__31539),
            .I(N__31501));
    Span4Mux_h I__6922 (
            .O(N__31534),
            .I(N__31501));
    Span4Mux_h I__6921 (
            .O(N__31531),
            .I(N__31498));
    Span4Mux_v I__6920 (
            .O(N__31528),
            .I(N__31493));
    Span4Mux_h I__6919 (
            .O(N__31525),
            .I(N__31493));
    Span4Mux_h I__6918 (
            .O(N__31520),
            .I(N__31488));
    Span4Mux_h I__6917 (
            .O(N__31517),
            .I(N__31488));
    Span4Mux_h I__6916 (
            .O(N__31512),
            .I(N__31483));
    LocalMux I__6915 (
            .O(N__31509),
            .I(N__31483));
    LocalMux I__6914 (
            .O(N__31506),
            .I(N__31480));
    Span4Mux_h I__6913 (
            .O(N__31501),
            .I(N__31477));
    Span4Mux_h I__6912 (
            .O(N__31498),
            .I(N__31474));
    Span4Mux_h I__6911 (
            .O(N__31493),
            .I(N__31469));
    Span4Mux_v I__6910 (
            .O(N__31488),
            .I(N__31469));
    Span4Mux_v I__6909 (
            .O(N__31483),
            .I(N__31464));
    Span4Mux_h I__6908 (
            .O(N__31480),
            .I(N__31464));
    Odrv4 I__6907 (
            .O(N__31477),
            .I(dataWriteZ0Z_2));
    Odrv4 I__6906 (
            .O(N__31474),
            .I(dataWriteZ0Z_2));
    Odrv4 I__6905 (
            .O(N__31469),
            .I(dataWriteZ0Z_2));
    Odrv4 I__6904 (
            .O(N__31464),
            .I(dataWriteZ0Z_2));
    CascadeMux I__6903 (
            .O(N__31455),
            .I(N__31452));
    InMux I__6902 (
            .O(N__31452),
            .I(N__31449));
    LocalMux I__6901 (
            .O(N__31449),
            .I(\PWMInstance2.PWMPulseWidthCountZ0Z_2 ));
    InMux I__6900 (
            .O(N__31446),
            .I(N__31443));
    LocalMux I__6899 (
            .O(N__31443),
            .I(OutReg_0_sqmuxa_0_a2_3_a2_2));
    CascadeMux I__6898 (
            .O(N__31440),
            .I(N__31431));
    CascadeMux I__6897 (
            .O(N__31439),
            .I(N__31426));
    CascadeMux I__6896 (
            .O(N__31438),
            .I(N__31423));
    InMux I__6895 (
            .O(N__31437),
            .I(N__31419));
    InMux I__6894 (
            .O(N__31436),
            .I(N__31416));
    InMux I__6893 (
            .O(N__31435),
            .I(N__31413));
    CascadeMux I__6892 (
            .O(N__31434),
            .I(N__31408));
    InMux I__6891 (
            .O(N__31431),
            .I(N__31404));
    InMux I__6890 (
            .O(N__31430),
            .I(N__31395));
    InMux I__6889 (
            .O(N__31429),
            .I(N__31395));
    InMux I__6888 (
            .O(N__31426),
            .I(N__31395));
    InMux I__6887 (
            .O(N__31423),
            .I(N__31395));
    InMux I__6886 (
            .O(N__31422),
            .I(N__31392));
    LocalMux I__6885 (
            .O(N__31419),
            .I(N__31389));
    LocalMux I__6884 (
            .O(N__31416),
            .I(N__31386));
    LocalMux I__6883 (
            .O(N__31413),
            .I(N__31383));
    InMux I__6882 (
            .O(N__31412),
            .I(N__31379));
    InMux I__6881 (
            .O(N__31411),
            .I(N__31375));
    InMux I__6880 (
            .O(N__31408),
            .I(N__31369));
    InMux I__6879 (
            .O(N__31407),
            .I(N__31369));
    LocalMux I__6878 (
            .O(N__31404),
            .I(N__31364));
    LocalMux I__6877 (
            .O(N__31395),
            .I(N__31364));
    LocalMux I__6876 (
            .O(N__31392),
            .I(N__31361));
    Span4Mux_v I__6875 (
            .O(N__31389),
            .I(N__31358));
    Span4Mux_v I__6874 (
            .O(N__31386),
            .I(N__31355));
    Span4Mux_v I__6873 (
            .O(N__31383),
            .I(N__31352));
    InMux I__6872 (
            .O(N__31382),
            .I(N__31349));
    LocalMux I__6871 (
            .O(N__31379),
            .I(N__31346));
    InMux I__6870 (
            .O(N__31378),
            .I(N__31343));
    LocalMux I__6869 (
            .O(N__31375),
            .I(N__31340));
    InMux I__6868 (
            .O(N__31374),
            .I(N__31337));
    LocalMux I__6867 (
            .O(N__31369),
            .I(N__31332));
    Span4Mux_h I__6866 (
            .O(N__31364),
            .I(N__31332));
    Span4Mux_v I__6865 (
            .O(N__31361),
            .I(N__31325));
    Span4Mux_h I__6864 (
            .O(N__31358),
            .I(N__31325));
    Span4Mux_h I__6863 (
            .O(N__31355),
            .I(N__31325));
    Span4Mux_v I__6862 (
            .O(N__31352),
            .I(N__31322));
    LocalMux I__6861 (
            .O(N__31349),
            .I(N__31317));
    Span4Mux_v I__6860 (
            .O(N__31346),
            .I(N__31317));
    LocalMux I__6859 (
            .O(N__31343),
            .I(N__31314));
    Span4Mux_h I__6858 (
            .O(N__31340),
            .I(N__31311));
    LocalMux I__6857 (
            .O(N__31337),
            .I(N__31308));
    Span4Mux_v I__6856 (
            .O(N__31332),
            .I(N__31303));
    Span4Mux_h I__6855 (
            .O(N__31325),
            .I(N__31303));
    Span4Mux_h I__6854 (
            .O(N__31322),
            .I(N__31298));
    Span4Mux_h I__6853 (
            .O(N__31317),
            .I(N__31298));
    Odrv12 I__6852 (
            .O(N__31314),
            .I(dataWriteZ0Z_0));
    Odrv4 I__6851 (
            .O(N__31311),
            .I(dataWriteZ0Z_0));
    Odrv12 I__6850 (
            .O(N__31308),
            .I(dataWriteZ0Z_0));
    Odrv4 I__6849 (
            .O(N__31303),
            .I(dataWriteZ0Z_0));
    Odrv4 I__6848 (
            .O(N__31298),
            .I(dataWriteZ0Z_0));
    InMux I__6847 (
            .O(N__31287),
            .I(N__31284));
    LocalMux I__6846 (
            .O(N__31284),
            .I(\PWMInstance2.PWMPulseWidthCountZ0Z_0 ));
    InMux I__6845 (
            .O(N__31281),
            .I(N__31275));
    InMux I__6844 (
            .O(N__31280),
            .I(N__31272));
    InMux I__6843 (
            .O(N__31279),
            .I(N__31268));
    InMux I__6842 (
            .O(N__31278),
            .I(N__31265));
    LocalMux I__6841 (
            .O(N__31275),
            .I(N__31261));
    LocalMux I__6840 (
            .O(N__31272),
            .I(N__31258));
    InMux I__6839 (
            .O(N__31271),
            .I(N__31253));
    LocalMux I__6838 (
            .O(N__31268),
            .I(N__31249));
    LocalMux I__6837 (
            .O(N__31265),
            .I(N__31244));
    InMux I__6836 (
            .O(N__31264),
            .I(N__31241));
    Span4Mux_v I__6835 (
            .O(N__31261),
            .I(N__31236));
    Span4Mux_v I__6834 (
            .O(N__31258),
            .I(N__31233));
    InMux I__6833 (
            .O(N__31257),
            .I(N__31230));
    InMux I__6832 (
            .O(N__31256),
            .I(N__31227));
    LocalMux I__6831 (
            .O(N__31253),
            .I(N__31224));
    InMux I__6830 (
            .O(N__31252),
            .I(N__31221));
    Span4Mux_h I__6829 (
            .O(N__31249),
            .I(N__31215));
    InMux I__6828 (
            .O(N__31248),
            .I(N__31212));
    InMux I__6827 (
            .O(N__31247),
            .I(N__31209));
    Span4Mux_v I__6826 (
            .O(N__31244),
            .I(N__31206));
    LocalMux I__6825 (
            .O(N__31241),
            .I(N__31203));
    InMux I__6824 (
            .O(N__31240),
            .I(N__31200));
    InMux I__6823 (
            .O(N__31239),
            .I(N__31197));
    Span4Mux_h I__6822 (
            .O(N__31236),
            .I(N__31190));
    Span4Mux_h I__6821 (
            .O(N__31233),
            .I(N__31190));
    LocalMux I__6820 (
            .O(N__31230),
            .I(N__31190));
    LocalMux I__6819 (
            .O(N__31227),
            .I(N__31187));
    Span4Mux_s2_v I__6818 (
            .O(N__31224),
            .I(N__31182));
    LocalMux I__6817 (
            .O(N__31221),
            .I(N__31182));
    InMux I__6816 (
            .O(N__31220),
            .I(N__31175));
    InMux I__6815 (
            .O(N__31219),
            .I(N__31175));
    InMux I__6814 (
            .O(N__31218),
            .I(N__31175));
    Span4Mux_v I__6813 (
            .O(N__31215),
            .I(N__31168));
    LocalMux I__6812 (
            .O(N__31212),
            .I(N__31168));
    LocalMux I__6811 (
            .O(N__31209),
            .I(N__31168));
    Span4Mux_h I__6810 (
            .O(N__31206),
            .I(N__31163));
    Span4Mux_v I__6809 (
            .O(N__31203),
            .I(N__31163));
    LocalMux I__6808 (
            .O(N__31200),
            .I(N__31158));
    LocalMux I__6807 (
            .O(N__31197),
            .I(N__31158));
    Span4Mux_v I__6806 (
            .O(N__31190),
            .I(N__31153));
    Span4Mux_h I__6805 (
            .O(N__31187),
            .I(N__31153));
    Span4Mux_v I__6804 (
            .O(N__31182),
            .I(N__31146));
    LocalMux I__6803 (
            .O(N__31175),
            .I(N__31146));
    Span4Mux_h I__6802 (
            .O(N__31168),
            .I(N__31146));
    Odrv4 I__6801 (
            .O(N__31163),
            .I(dataWriteZ0Z_1));
    Odrv12 I__6800 (
            .O(N__31158),
            .I(dataWriteZ0Z_1));
    Odrv4 I__6799 (
            .O(N__31153),
            .I(dataWriteZ0Z_1));
    Odrv4 I__6798 (
            .O(N__31146),
            .I(dataWriteZ0Z_1));
    InMux I__6797 (
            .O(N__31137),
            .I(N__31134));
    LocalMux I__6796 (
            .O(N__31134),
            .I(\PWMInstance2.PWMPulseWidthCountZ0Z_1 ));
    InMux I__6795 (
            .O(N__31131),
            .I(N__31128));
    LocalMux I__6794 (
            .O(N__31128),
            .I(\PWMInstance2.PWMPulseWidthCountZ0Z_7 ));
    InMux I__6793 (
            .O(N__31125),
            .I(N__31121));
    InMux I__6792 (
            .O(N__31124),
            .I(N__31115));
    LocalMux I__6791 (
            .O(N__31121),
            .I(N__31104));
    InMux I__6790 (
            .O(N__31120),
            .I(N__31101));
    InMux I__6789 (
            .O(N__31119),
            .I(N__31098));
    InMux I__6788 (
            .O(N__31118),
            .I(N__31095));
    LocalMux I__6787 (
            .O(N__31115),
            .I(N__31091));
    InMux I__6786 (
            .O(N__31114),
            .I(N__31088));
    InMux I__6785 (
            .O(N__31113),
            .I(N__31082));
    InMux I__6784 (
            .O(N__31112),
            .I(N__31082));
    InMux I__6783 (
            .O(N__31111),
            .I(N__31079));
    InMux I__6782 (
            .O(N__31110),
            .I(N__31076));
    InMux I__6781 (
            .O(N__31109),
            .I(N__31073));
    InMux I__6780 (
            .O(N__31108),
            .I(N__31070));
    InMux I__6779 (
            .O(N__31107),
            .I(N__31067));
    Span4Mux_v I__6778 (
            .O(N__31104),
            .I(N__31064));
    LocalMux I__6777 (
            .O(N__31101),
            .I(N__31060));
    LocalMux I__6776 (
            .O(N__31098),
            .I(N__31057));
    LocalMux I__6775 (
            .O(N__31095),
            .I(N__31054));
    InMux I__6774 (
            .O(N__31094),
            .I(N__31051));
    Span4Mux_v I__6773 (
            .O(N__31091),
            .I(N__31048));
    LocalMux I__6772 (
            .O(N__31088),
            .I(N__31045));
    InMux I__6771 (
            .O(N__31087),
            .I(N__31042));
    LocalMux I__6770 (
            .O(N__31082),
            .I(N__31037));
    LocalMux I__6769 (
            .O(N__31079),
            .I(N__31037));
    LocalMux I__6768 (
            .O(N__31076),
            .I(N__31032));
    LocalMux I__6767 (
            .O(N__31073),
            .I(N__31032));
    LocalMux I__6766 (
            .O(N__31070),
            .I(N__31027));
    LocalMux I__6765 (
            .O(N__31067),
            .I(N__31027));
    Span4Mux_h I__6764 (
            .O(N__31064),
            .I(N__31024));
    InMux I__6763 (
            .O(N__31063),
            .I(N__31021));
    Span4Mux_v I__6762 (
            .O(N__31060),
            .I(N__31018));
    Span4Mux_h I__6761 (
            .O(N__31057),
            .I(N__31011));
    Span4Mux_v I__6760 (
            .O(N__31054),
            .I(N__31011));
    LocalMux I__6759 (
            .O(N__31051),
            .I(N__31011));
    Span4Mux_v I__6758 (
            .O(N__31048),
            .I(N__31004));
    Span4Mux_v I__6757 (
            .O(N__31045),
            .I(N__31004));
    LocalMux I__6756 (
            .O(N__31042),
            .I(N__31004));
    Span4Mux_v I__6755 (
            .O(N__31037),
            .I(N__31001));
    Span4Mux_h I__6754 (
            .O(N__31032),
            .I(N__30996));
    Span4Mux_h I__6753 (
            .O(N__31027),
            .I(N__30996));
    Span4Mux_h I__6752 (
            .O(N__31024),
            .I(N__30991));
    LocalMux I__6751 (
            .O(N__31021),
            .I(N__30991));
    Span4Mux_v I__6750 (
            .O(N__31018),
            .I(N__30988));
    Span4Mux_v I__6749 (
            .O(N__31011),
            .I(N__30981));
    Span4Mux_h I__6748 (
            .O(N__31004),
            .I(N__30981));
    Span4Mux_v I__6747 (
            .O(N__31001),
            .I(N__30981));
    Span4Mux_v I__6746 (
            .O(N__30996),
            .I(N__30978));
    Odrv4 I__6745 (
            .O(N__30991),
            .I(dataWriteZ0Z_6));
    Odrv4 I__6744 (
            .O(N__30988),
            .I(dataWriteZ0Z_6));
    Odrv4 I__6743 (
            .O(N__30981),
            .I(dataWriteZ0Z_6));
    Odrv4 I__6742 (
            .O(N__30978),
            .I(dataWriteZ0Z_6));
    InMux I__6741 (
            .O(N__30969),
            .I(N__30966));
    LocalMux I__6740 (
            .O(N__30966),
            .I(\PWMInstance2.PWMPulseWidthCountZ0Z_6 ));
    InMux I__6739 (
            .O(N__30963),
            .I(N__30960));
    LocalMux I__6738 (
            .O(N__30960),
            .I(\PWMInstance2.PWMPulseWidthCountZ0Z_8 ));
    InMux I__6737 (
            .O(N__30957),
            .I(N__30954));
    LocalMux I__6736 (
            .O(N__30954),
            .I(\PWMInstance2.PWMPulseWidthCountZ0Z_9 ));
    InMux I__6735 (
            .O(N__30951),
            .I(N__30948));
    LocalMux I__6734 (
            .O(N__30948),
            .I(N__30944));
    CascadeMux I__6733 (
            .O(N__30947),
            .I(N__30940));
    Span4Mux_h I__6732 (
            .O(N__30944),
            .I(N__30937));
    CascadeMux I__6731 (
            .O(N__30943),
            .I(N__30934));
    InMux I__6730 (
            .O(N__30940),
            .I(N__30931));
    Span4Mux_h I__6729 (
            .O(N__30937),
            .I(N__30928));
    InMux I__6728 (
            .O(N__30934),
            .I(N__30925));
    LocalMux I__6727 (
            .O(N__30931),
            .I(dataRead1_0));
    Odrv4 I__6726 (
            .O(N__30928),
            .I(dataRead1_0));
    LocalMux I__6725 (
            .O(N__30925),
            .I(dataRead1_0));
    CascadeMux I__6724 (
            .O(N__30918),
            .I(OutReg_0_5_i_m3_ns_1_0_cascade_));
    InMux I__6723 (
            .O(N__30915),
            .I(N__30912));
    LocalMux I__6722 (
            .O(N__30912),
            .I(N__30909));
    Span4Mux_h I__6721 (
            .O(N__30909),
            .I(N__30904));
    CascadeMux I__6720 (
            .O(N__30908),
            .I(N__30901));
    InMux I__6719 (
            .O(N__30907),
            .I(N__30898));
    Span4Mux_v I__6718 (
            .O(N__30904),
            .I(N__30895));
    InMux I__6717 (
            .O(N__30901),
            .I(N__30892));
    LocalMux I__6716 (
            .O(N__30898),
            .I(dataRead5_0));
    Odrv4 I__6715 (
            .O(N__30895),
            .I(dataRead5_0));
    LocalMux I__6714 (
            .O(N__30892),
            .I(dataRead5_0));
    CascadeMux I__6713 (
            .O(N__30885),
            .I(OutReg_ess_RNO_1Z0Z_0_cascade_));
    InMux I__6712 (
            .O(N__30882),
            .I(N__30879));
    LocalMux I__6711 (
            .O(N__30879),
            .I(N__30874));
    CascadeMux I__6710 (
            .O(N__30878),
            .I(N__30871));
    InMux I__6709 (
            .O(N__30877),
            .I(N__30868));
    Span4Mux_v I__6708 (
            .O(N__30874),
            .I(N__30865));
    InMux I__6707 (
            .O(N__30871),
            .I(N__30862));
    LocalMux I__6706 (
            .O(N__30868),
            .I(N__30857));
    Span4Mux_h I__6705 (
            .O(N__30865),
            .I(N__30857));
    LocalMux I__6704 (
            .O(N__30862),
            .I(N__30854));
    Odrv4 I__6703 (
            .O(N__30857),
            .I(dataRead3_0));
    Odrv12 I__6702 (
            .O(N__30854),
            .I(dataRead3_0));
    CascadeMux I__6701 (
            .O(N__30849),
            .I(N__30846));
    InMux I__6700 (
            .O(N__30846),
            .I(N__30842));
    CascadeMux I__6699 (
            .O(N__30845),
            .I(N__30839));
    LocalMux I__6698 (
            .O(N__30842),
            .I(N__30835));
    InMux I__6697 (
            .O(N__30839),
            .I(N__30832));
    InMux I__6696 (
            .O(N__30838),
            .I(N__30829));
    Span4Mux_v I__6695 (
            .O(N__30835),
            .I(N__30826));
    LocalMux I__6694 (
            .O(N__30832),
            .I(N__30823));
    LocalMux I__6693 (
            .O(N__30829),
            .I(N__30818));
    Span4Mux_h I__6692 (
            .O(N__30826),
            .I(N__30818));
    Span4Mux_h I__6691 (
            .O(N__30823),
            .I(N__30815));
    Odrv4 I__6690 (
            .O(N__30818),
            .I(dataRead2_0));
    Odrv4 I__6689 (
            .O(N__30815),
            .I(dataRead2_0));
    CascadeMux I__6688 (
            .O(N__30810),
            .I(N__30806));
    InMux I__6687 (
            .O(N__30809),
            .I(N__30803));
    InMux I__6686 (
            .O(N__30806),
            .I(N__30800));
    LocalMux I__6685 (
            .O(N__30803),
            .I(N__30796));
    LocalMux I__6684 (
            .O(N__30800),
            .I(N__30793));
    InMux I__6683 (
            .O(N__30799),
            .I(N__30790));
    Span4Mux_h I__6682 (
            .O(N__30796),
            .I(N__30785));
    Span4Mux_h I__6681 (
            .O(N__30793),
            .I(N__30785));
    LocalMux I__6680 (
            .O(N__30790),
            .I(dataRead6_0));
    Odrv4 I__6679 (
            .O(N__30785),
            .I(dataRead6_0));
    CascadeMux I__6678 (
            .O(N__30780),
            .I(OutReg_0_4_i_m3_ns_1_0_cascade_));
    InMux I__6677 (
            .O(N__30777),
            .I(N__30773));
    CascadeMux I__6676 (
            .O(N__30776),
            .I(N__30770));
    LocalMux I__6675 (
            .O(N__30773),
            .I(N__30766));
    InMux I__6674 (
            .O(N__30770),
            .I(N__30763));
    InMux I__6673 (
            .O(N__30769),
            .I(N__30760));
    Span4Mux_h I__6672 (
            .O(N__30766),
            .I(N__30757));
    LocalMux I__6671 (
            .O(N__30763),
            .I(N__30754));
    LocalMux I__6670 (
            .O(N__30760),
            .I(dataRead7_0));
    Odrv4 I__6669 (
            .O(N__30757),
            .I(dataRead7_0));
    Odrv12 I__6668 (
            .O(N__30754),
            .I(dataRead7_0));
    InMux I__6667 (
            .O(N__30747),
            .I(N__30744));
    LocalMux I__6666 (
            .O(N__30744),
            .I(OutReg_ess_RNO_0Z0Z_0));
    CascadeMux I__6665 (
            .O(N__30741),
            .I(N__30738));
    InMux I__6664 (
            .O(N__30738),
            .I(N__30735));
    LocalMux I__6663 (
            .O(N__30735),
            .I(N__30732));
    Odrv4 I__6662 (
            .O(N__30732),
            .I(OutRegZ0Z_0));
    InMux I__6661 (
            .O(N__30729),
            .I(N__30726));
    LocalMux I__6660 (
            .O(N__30726),
            .I(N__30723));
    Span4Mux_h I__6659 (
            .O(N__30723),
            .I(N__30720));
    Odrv4 I__6658 (
            .O(N__30720),
            .I(OutReg_ess_RNO_0Z0Z_1));
    InMux I__6657 (
            .O(N__30717),
            .I(N__30714));
    LocalMux I__6656 (
            .O(N__30714),
            .I(OutRegZ0Z_1));
    InMux I__6655 (
            .O(N__30711),
            .I(N__30707));
    InMux I__6654 (
            .O(N__30710),
            .I(N__30704));
    LocalMux I__6653 (
            .O(N__30707),
            .I(N__30700));
    LocalMux I__6652 (
            .O(N__30704),
            .I(N__30697));
    InMux I__6651 (
            .O(N__30703),
            .I(N__30694));
    Span4Mux_v I__6650 (
            .O(N__30700),
            .I(N__30691));
    Span4Mux_h I__6649 (
            .O(N__30697),
            .I(N__30688));
    LocalMux I__6648 (
            .O(N__30694),
            .I(N__30685));
    Span4Mux_h I__6647 (
            .O(N__30691),
            .I(N__30680));
    Span4Mux_h I__6646 (
            .O(N__30688),
            .I(N__30680));
    Odrv12 I__6645 (
            .O(N__30685),
            .I(dataRead2_8));
    Odrv4 I__6644 (
            .O(N__30680),
            .I(dataRead2_8));
    CascadeMux I__6643 (
            .O(N__30675),
            .I(N__30672));
    InMux I__6642 (
            .O(N__30672),
            .I(N__30669));
    LocalMux I__6641 (
            .O(N__30669),
            .I(N__30665));
    InMux I__6640 (
            .O(N__30668),
            .I(N__30662));
    Span4Mux_h I__6639 (
            .O(N__30665),
            .I(N__30658));
    LocalMux I__6638 (
            .O(N__30662),
            .I(N__30655));
    InMux I__6637 (
            .O(N__30661),
            .I(N__30652));
    Span4Mux_h I__6636 (
            .O(N__30658),
            .I(N__30649));
    Odrv4 I__6635 (
            .O(N__30655),
            .I(dataRead3_8));
    LocalMux I__6634 (
            .O(N__30652),
            .I(dataRead3_8));
    Odrv4 I__6633 (
            .O(N__30649),
            .I(dataRead3_8));
    CascadeMux I__6632 (
            .O(N__30642),
            .I(N__30639));
    InMux I__6631 (
            .O(N__30639),
            .I(N__30635));
    InMux I__6630 (
            .O(N__30638),
            .I(N__30631));
    LocalMux I__6629 (
            .O(N__30635),
            .I(N__30628));
    InMux I__6628 (
            .O(N__30634),
            .I(N__30625));
    LocalMux I__6627 (
            .O(N__30631),
            .I(N__30622));
    Span4Mux_h I__6626 (
            .O(N__30628),
            .I(N__30616));
    LocalMux I__6625 (
            .O(N__30625),
            .I(N__30616));
    Span4Mux_h I__6624 (
            .O(N__30622),
            .I(N__30613));
    InMux I__6623 (
            .O(N__30621),
            .I(N__30610));
    Span4Mux_h I__6622 (
            .O(N__30616),
            .I(N__30607));
    Odrv4 I__6621 (
            .O(N__30613),
            .I(data_receivedZ0Z_3));
    LocalMux I__6620 (
            .O(N__30610),
            .I(data_receivedZ0Z_3));
    Odrv4 I__6619 (
            .O(N__30607),
            .I(data_receivedZ0Z_3));
    CascadeMux I__6618 (
            .O(N__30600),
            .I(data_received_esr_RNI7L871Z0Z_3_cascade_));
    InMux I__6617 (
            .O(N__30597),
            .I(\QuadInstance0.un1_Quad_cry_13 ));
    InMux I__6616 (
            .O(N__30594),
            .I(N__30591));
    LocalMux I__6615 (
            .O(N__30591),
            .I(N__30588));
    Odrv4 I__6614 (
            .O(N__30588),
            .I(\QuadInstance0.un1_Quad_axb_15 ));
    InMux I__6613 (
            .O(N__30585),
            .I(\QuadInstance0.un1_Quad_cry_14 ));
    InMux I__6612 (
            .O(N__30582),
            .I(N__30576));
    InMux I__6611 (
            .O(N__30581),
            .I(N__30576));
    LocalMux I__6610 (
            .O(N__30576),
            .I(N__30573));
    Odrv4 I__6609 (
            .O(N__30573),
            .I(dataRead0_15));
    InMux I__6608 (
            .O(N__30570),
            .I(N__30565));
    InMux I__6607 (
            .O(N__30569),
            .I(N__30562));
    InMux I__6606 (
            .O(N__30568),
            .I(N__30559));
    LocalMux I__6605 (
            .O(N__30565),
            .I(N__30556));
    LocalMux I__6604 (
            .O(N__30562),
            .I(N__30551));
    LocalMux I__6603 (
            .O(N__30559),
            .I(N__30551));
    Span4Mux_v I__6602 (
            .O(N__30556),
            .I(N__30548));
    Span4Mux_h I__6601 (
            .O(N__30551),
            .I(N__30545));
    Sp12to4 I__6600 (
            .O(N__30548),
            .I(N__30542));
    Span4Mux_h I__6599 (
            .O(N__30545),
            .I(N__30539));
    Odrv12 I__6598 (
            .O(N__30542),
            .I(dataRead1_2));
    Odrv4 I__6597 (
            .O(N__30539),
            .I(dataRead1_2));
    CascadeMux I__6596 (
            .O(N__30534),
            .I(N__30531));
    InMux I__6595 (
            .O(N__30531),
            .I(N__30527));
    InMux I__6594 (
            .O(N__30530),
            .I(N__30523));
    LocalMux I__6593 (
            .O(N__30527),
            .I(N__30520));
    InMux I__6592 (
            .O(N__30526),
            .I(N__30517));
    LocalMux I__6591 (
            .O(N__30523),
            .I(N__30514));
    Span4Mux_h I__6590 (
            .O(N__30520),
            .I(N__30511));
    LocalMux I__6589 (
            .O(N__30517),
            .I(N__30508));
    Span4Mux_h I__6588 (
            .O(N__30514),
            .I(N__30505));
    Span4Mux_h I__6587 (
            .O(N__30511),
            .I(N__30502));
    Span4Mux_v I__6586 (
            .O(N__30508),
            .I(N__30499));
    Odrv4 I__6585 (
            .O(N__30505),
            .I(dataRead5_2));
    Odrv4 I__6584 (
            .O(N__30502),
            .I(dataRead5_2));
    Odrv4 I__6583 (
            .O(N__30499),
            .I(dataRead5_2));
    InMux I__6582 (
            .O(N__30492),
            .I(N__30489));
    LocalMux I__6581 (
            .O(N__30489),
            .I(N__30486));
    Span4Mux_v I__6580 (
            .O(N__30486),
            .I(N__30483));
    Odrv4 I__6579 (
            .O(N__30483),
            .I(OutReg_0_5_i_m3_ns_1_2));
    CascadeMux I__6578 (
            .O(N__30480),
            .I(OutReg_esr_RNO_2Z0Z_2_cascade_));
    CascadeMux I__6577 (
            .O(N__30477),
            .I(OutReg_esr_RNO_0Z0Z_2_cascade_));
    InMux I__6576 (
            .O(N__30474),
            .I(N__30471));
    LocalMux I__6575 (
            .O(N__30471),
            .I(N__30468));
    Odrv4 I__6574 (
            .O(N__30468),
            .I(OutRegZ0Z_2));
    InMux I__6573 (
            .O(N__30465),
            .I(N__30462));
    LocalMux I__6572 (
            .O(N__30462),
            .I(N__30457));
    InMux I__6571 (
            .O(N__30461),
            .I(N__30454));
    InMux I__6570 (
            .O(N__30460),
            .I(N__30451));
    Span4Mux_v I__6569 (
            .O(N__30457),
            .I(N__30446));
    LocalMux I__6568 (
            .O(N__30454),
            .I(N__30446));
    LocalMux I__6567 (
            .O(N__30451),
            .I(N__30443));
    Span4Mux_h I__6566 (
            .O(N__30446),
            .I(N__30440));
    Span4Mux_v I__6565 (
            .O(N__30443),
            .I(N__30437));
    Span4Mux_h I__6564 (
            .O(N__30440),
            .I(N__30434));
    Span4Mux_h I__6563 (
            .O(N__30437),
            .I(N__30431));
    Odrv4 I__6562 (
            .O(N__30434),
            .I(dataRead2_2));
    Odrv4 I__6561 (
            .O(N__30431),
            .I(dataRead2_2));
    CascadeMux I__6560 (
            .O(N__30426),
            .I(N__30423));
    InMux I__6559 (
            .O(N__30423),
            .I(N__30419));
    InMux I__6558 (
            .O(N__30422),
            .I(N__30415));
    LocalMux I__6557 (
            .O(N__30419),
            .I(N__30412));
    InMux I__6556 (
            .O(N__30418),
            .I(N__30409));
    LocalMux I__6555 (
            .O(N__30415),
            .I(N__30406));
    Span4Mux_h I__6554 (
            .O(N__30412),
            .I(N__30403));
    LocalMux I__6553 (
            .O(N__30409),
            .I(N__30400));
    Sp12to4 I__6552 (
            .O(N__30406),
            .I(N__30397));
    Span4Mux_v I__6551 (
            .O(N__30403),
            .I(N__30392));
    Span4Mux_v I__6550 (
            .O(N__30400),
            .I(N__30392));
    Odrv12 I__6549 (
            .O(N__30397),
            .I(dataRead3_2));
    Odrv4 I__6548 (
            .O(N__30392),
            .I(dataRead3_2));
    InMux I__6547 (
            .O(N__30387),
            .I(N__30383));
    InMux I__6546 (
            .O(N__30386),
            .I(N__30380));
    LocalMux I__6545 (
            .O(N__30383),
            .I(N__30376));
    LocalMux I__6544 (
            .O(N__30380),
            .I(N__30373));
    InMux I__6543 (
            .O(N__30379),
            .I(N__30370));
    Span4Mux_v I__6542 (
            .O(N__30376),
            .I(N__30367));
    Span4Mux_v I__6541 (
            .O(N__30373),
            .I(N__30362));
    LocalMux I__6540 (
            .O(N__30370),
            .I(N__30362));
    Span4Mux_h I__6539 (
            .O(N__30367),
            .I(N__30357));
    Span4Mux_v I__6538 (
            .O(N__30362),
            .I(N__30357));
    Odrv4 I__6537 (
            .O(N__30357),
            .I(dataRead7_2));
    InMux I__6536 (
            .O(N__30354),
            .I(N__30350));
    InMux I__6535 (
            .O(N__30353),
            .I(N__30347));
    LocalMux I__6534 (
            .O(N__30350),
            .I(N__30341));
    LocalMux I__6533 (
            .O(N__30347),
            .I(N__30341));
    InMux I__6532 (
            .O(N__30346),
            .I(N__30338));
    Span12Mux_h I__6531 (
            .O(N__30341),
            .I(N__30335));
    LocalMux I__6530 (
            .O(N__30338),
            .I(N__30332));
    Odrv12 I__6529 (
            .O(N__30335),
            .I(dataRead6_2));
    Odrv4 I__6528 (
            .O(N__30332),
            .I(dataRead6_2));
    CascadeMux I__6527 (
            .O(N__30327),
            .I(OutReg_0_4_i_m3_ns_1_2_cascade_));
    InMux I__6526 (
            .O(N__30324),
            .I(N__30321));
    LocalMux I__6525 (
            .O(N__30321),
            .I(OutReg_esr_RNO_1Z0Z_2));
    InMux I__6524 (
            .O(N__30318),
            .I(N__30314));
    CascadeMux I__6523 (
            .O(N__30317),
            .I(N__30311));
    LocalMux I__6522 (
            .O(N__30314),
            .I(N__30308));
    InMux I__6521 (
            .O(N__30311),
            .I(N__30305));
    Span4Mux_v I__6520 (
            .O(N__30308),
            .I(N__30300));
    LocalMux I__6519 (
            .O(N__30305),
            .I(N__30300));
    Span4Mux_h I__6518 (
            .O(N__30300),
            .I(N__30296));
    InMux I__6517 (
            .O(N__30299),
            .I(N__30293));
    Span4Mux_h I__6516 (
            .O(N__30296),
            .I(N__30290));
    LocalMux I__6515 (
            .O(N__30293),
            .I(dataRead0_0));
    Odrv4 I__6514 (
            .O(N__30290),
            .I(dataRead0_0));
    CascadeMux I__6513 (
            .O(N__30285),
            .I(N__30281));
    CascadeMux I__6512 (
            .O(N__30284),
            .I(N__30278));
    InMux I__6511 (
            .O(N__30281),
            .I(N__30275));
    InMux I__6510 (
            .O(N__30278),
            .I(N__30272));
    LocalMux I__6509 (
            .O(N__30275),
            .I(N__30269));
    LocalMux I__6508 (
            .O(N__30272),
            .I(N__30265));
    Span4Mux_v I__6507 (
            .O(N__30269),
            .I(N__30262));
    InMux I__6506 (
            .O(N__30268),
            .I(N__30259));
    Span4Mux_s2_v I__6505 (
            .O(N__30265),
            .I(N__30256));
    Span4Mux_h I__6504 (
            .O(N__30262),
            .I(N__30253));
    LocalMux I__6503 (
            .O(N__30259),
            .I(N__30248));
    Span4Mux_h I__6502 (
            .O(N__30256),
            .I(N__30248));
    Odrv4 I__6501 (
            .O(N__30253),
            .I(dataRead4_0));
    Odrv4 I__6500 (
            .O(N__30248),
            .I(dataRead4_0));
    InMux I__6499 (
            .O(N__30243),
            .I(N__30240));
    LocalMux I__6498 (
            .O(N__30240),
            .I(N__30237));
    Span4Mux_h I__6497 (
            .O(N__30237),
            .I(N__30234));
    Odrv4 I__6496 (
            .O(N__30234),
            .I(\QuadInstance0.Quad_RNO_0_0_6 ));
    InMux I__6495 (
            .O(N__30231),
            .I(\QuadInstance0.un1_Quad_cry_5 ));
    InMux I__6494 (
            .O(N__30228),
            .I(N__30223));
    InMux I__6493 (
            .O(N__30227),
            .I(N__30218));
    InMux I__6492 (
            .O(N__30226),
            .I(N__30218));
    LocalMux I__6491 (
            .O(N__30223),
            .I(dataRead0_7));
    LocalMux I__6490 (
            .O(N__30218),
            .I(dataRead0_7));
    CascadeMux I__6489 (
            .O(N__30213),
            .I(N__30210));
    InMux I__6488 (
            .O(N__30210),
            .I(N__30207));
    LocalMux I__6487 (
            .O(N__30207),
            .I(\QuadInstance0.Quad_RNIMKBH1Z0Z_7 ));
    InMux I__6486 (
            .O(N__30204),
            .I(N__30201));
    LocalMux I__6485 (
            .O(N__30201),
            .I(\QuadInstance0.Quad_RNO_0_0_7 ));
    InMux I__6484 (
            .O(N__30198),
            .I(\QuadInstance0.un1_Quad_cry_6 ));
    InMux I__6483 (
            .O(N__30195),
            .I(N__30190));
    InMux I__6482 (
            .O(N__30194),
            .I(N__30185));
    InMux I__6481 (
            .O(N__30193),
            .I(N__30185));
    LocalMux I__6480 (
            .O(N__30190),
            .I(dataRead0_8));
    LocalMux I__6479 (
            .O(N__30185),
            .I(dataRead0_8));
    CascadeMux I__6478 (
            .O(N__30180),
            .I(N__30177));
    InMux I__6477 (
            .O(N__30177),
            .I(N__30174));
    LocalMux I__6476 (
            .O(N__30174),
            .I(\QuadInstance0.Quad_RNINLBH1Z0Z_8 ));
    InMux I__6475 (
            .O(N__30171),
            .I(N__30168));
    LocalMux I__6474 (
            .O(N__30168),
            .I(\QuadInstance0.Quad_RNO_0_0_8 ));
    InMux I__6473 (
            .O(N__30165),
            .I(bfn_17_7_0_));
    InMux I__6472 (
            .O(N__30162),
            .I(N__30158));
    InMux I__6471 (
            .O(N__30161),
            .I(N__30154));
    LocalMux I__6470 (
            .O(N__30158),
            .I(N__30151));
    InMux I__6469 (
            .O(N__30157),
            .I(N__30148));
    LocalMux I__6468 (
            .O(N__30154),
            .I(N__30145));
    Span4Mux_v I__6467 (
            .O(N__30151),
            .I(N__30140));
    LocalMux I__6466 (
            .O(N__30148),
            .I(N__30140));
    Span4Mux_v I__6465 (
            .O(N__30145),
            .I(N__30137));
    Span4Mux_h I__6464 (
            .O(N__30140),
            .I(N__30134));
    Odrv4 I__6463 (
            .O(N__30137),
            .I(dataRead0_9));
    Odrv4 I__6462 (
            .O(N__30134),
            .I(dataRead0_9));
    CascadeMux I__6461 (
            .O(N__30129),
            .I(N__30126));
    InMux I__6460 (
            .O(N__30126),
            .I(N__30123));
    LocalMux I__6459 (
            .O(N__30123),
            .I(N__30120));
    Odrv4 I__6458 (
            .O(N__30120),
            .I(\QuadInstance0.Quad_RNIOMBH1Z0Z_9 ));
    InMux I__6457 (
            .O(N__30117),
            .I(N__30114));
    LocalMux I__6456 (
            .O(N__30114),
            .I(N__30111));
    Span4Mux_h I__6455 (
            .O(N__30111),
            .I(N__30108));
    Odrv4 I__6454 (
            .O(N__30108),
            .I(\QuadInstance0.Quad_RNO_0_0_9 ));
    InMux I__6453 (
            .O(N__30105),
            .I(\QuadInstance0.un1_Quad_cry_8 ));
    InMux I__6452 (
            .O(N__30102),
            .I(\QuadInstance0.un1_Quad_cry_9 ));
    InMux I__6451 (
            .O(N__30099),
            .I(N__30094));
    InMux I__6450 (
            .O(N__30098),
            .I(N__30091));
    InMux I__6449 (
            .O(N__30097),
            .I(N__30088));
    LocalMux I__6448 (
            .O(N__30094),
            .I(N__30083));
    LocalMux I__6447 (
            .O(N__30091),
            .I(N__30083));
    LocalMux I__6446 (
            .O(N__30088),
            .I(N__30080));
    Odrv12 I__6445 (
            .O(N__30083),
            .I(dataRead0_11));
    Odrv12 I__6444 (
            .O(N__30080),
            .I(dataRead0_11));
    CascadeMux I__6443 (
            .O(N__30075),
            .I(N__30072));
    InMux I__6442 (
            .O(N__30072),
            .I(N__30069));
    LocalMux I__6441 (
            .O(N__30069),
            .I(\QuadInstance0.Quad_RNI1M8Q1Z0Z_11 ));
    InMux I__6440 (
            .O(N__30066),
            .I(N__30063));
    LocalMux I__6439 (
            .O(N__30063),
            .I(N__30060));
    Odrv12 I__6438 (
            .O(N__30060),
            .I(\QuadInstance0.Quad_RNO_0_0_11 ));
    InMux I__6437 (
            .O(N__30057),
            .I(\QuadInstance0.un1_Quad_cry_10 ));
    InMux I__6436 (
            .O(N__30054),
            .I(N__30050));
    InMux I__6435 (
            .O(N__30053),
            .I(N__30046));
    LocalMux I__6434 (
            .O(N__30050),
            .I(N__30043));
    InMux I__6433 (
            .O(N__30049),
            .I(N__30040));
    LocalMux I__6432 (
            .O(N__30046),
            .I(dataRead0_12));
    Odrv4 I__6431 (
            .O(N__30043),
            .I(dataRead0_12));
    LocalMux I__6430 (
            .O(N__30040),
            .I(dataRead0_12));
    CascadeMux I__6429 (
            .O(N__30033),
            .I(N__30030));
    InMux I__6428 (
            .O(N__30030),
            .I(N__30027));
    LocalMux I__6427 (
            .O(N__30027),
            .I(\QuadInstance0.Quad_RNI2N8Q1Z0Z_12 ));
    InMux I__6426 (
            .O(N__30024),
            .I(N__30021));
    LocalMux I__6425 (
            .O(N__30021),
            .I(\QuadInstance0.Quad_RNO_0_0_12 ));
    InMux I__6424 (
            .O(N__30018),
            .I(\QuadInstance0.un1_Quad_cry_11 ));
    CascadeMux I__6423 (
            .O(N__30015),
            .I(N__30010));
    InMux I__6422 (
            .O(N__30014),
            .I(N__30007));
    InMux I__6421 (
            .O(N__30013),
            .I(N__30002));
    InMux I__6420 (
            .O(N__30010),
            .I(N__30002));
    LocalMux I__6419 (
            .O(N__30007),
            .I(dataRead0_13));
    LocalMux I__6418 (
            .O(N__30002),
            .I(dataRead0_13));
    CascadeMux I__6417 (
            .O(N__29997),
            .I(N__29994));
    InMux I__6416 (
            .O(N__29994),
            .I(N__29991));
    LocalMux I__6415 (
            .O(N__29991),
            .I(\QuadInstance0.Quad_RNI3O8Q1Z0Z_13 ));
    InMux I__6414 (
            .O(N__29988),
            .I(N__29985));
    LocalMux I__6413 (
            .O(N__29985),
            .I(\QuadInstance0.Quad_RNO_0_0_13 ));
    InMux I__6412 (
            .O(N__29982),
            .I(\QuadInstance0.un1_Quad_cry_12 ));
    InMux I__6411 (
            .O(N__29979),
            .I(N__29976));
    LocalMux I__6410 (
            .O(N__29976),
            .I(N__29973));
    Odrv4 I__6409 (
            .O(N__29973),
            .I(\QuadInstance4.Quad_RNO_0_4_14 ));
    CascadeMux I__6408 (
            .O(N__29970),
            .I(N__29966));
    CascadeMux I__6407 (
            .O(N__29969),
            .I(N__29962));
    InMux I__6406 (
            .O(N__29966),
            .I(N__29959));
    CascadeMux I__6405 (
            .O(N__29965),
            .I(N__29956));
    InMux I__6404 (
            .O(N__29962),
            .I(N__29953));
    LocalMux I__6403 (
            .O(N__29959),
            .I(N__29950));
    InMux I__6402 (
            .O(N__29956),
            .I(N__29947));
    LocalMux I__6401 (
            .O(N__29953),
            .I(N__29944));
    Span4Mux_v I__6400 (
            .O(N__29950),
            .I(N__29941));
    LocalMux I__6399 (
            .O(N__29947),
            .I(dataRead4_14));
    Odrv12 I__6398 (
            .O(N__29944),
            .I(dataRead4_14));
    Odrv4 I__6397 (
            .O(N__29941),
            .I(dataRead4_14));
    InMux I__6396 (
            .O(N__29934),
            .I(N__29931));
    LocalMux I__6395 (
            .O(N__29931),
            .I(N__29928));
    Span4Mux_v I__6394 (
            .O(N__29928),
            .I(N__29925));
    Sp12to4 I__6393 (
            .O(N__29925),
            .I(N__29922));
    Odrv12 I__6392 (
            .O(N__29922),
            .I(\QuadInstance0.delayedCh_BZ0Z_0 ));
    InMux I__6391 (
            .O(N__29919),
            .I(N__29916));
    LocalMux I__6390 (
            .O(N__29916),
            .I(N__29913));
    Span4Mux_h I__6389 (
            .O(N__29913),
            .I(N__29910));
    Odrv4 I__6388 (
            .O(N__29910),
            .I(\QuadInstance4.delayedCh_BZ0Z_0 ));
    CascadeMux I__6387 (
            .O(N__29907),
            .I(N__29903));
    InMux I__6386 (
            .O(N__29906),
            .I(N__29900));
    InMux I__6385 (
            .O(N__29903),
            .I(N__29897));
    LocalMux I__6384 (
            .O(N__29900),
            .I(\QuadInstance4.delayedCh_BZ0Z_1 ));
    LocalMux I__6383 (
            .O(N__29897),
            .I(\QuadInstance4.delayedCh_BZ0Z_1 ));
    InMux I__6382 (
            .O(N__29892),
            .I(N__29889));
    LocalMux I__6381 (
            .O(N__29889),
            .I(N__29886));
    Span4Mux_h I__6380 (
            .O(N__29886),
            .I(N__29883));
    Odrv4 I__6379 (
            .O(N__29883),
            .I(\QuadInstance0.Quad_RNO_0Z0Z_1 ));
    InMux I__6378 (
            .O(N__29880),
            .I(\QuadInstance0.un1_Quad_cry_0 ));
    InMux I__6377 (
            .O(N__29877),
            .I(N__29874));
    LocalMux I__6376 (
            .O(N__29874),
            .I(N__29871));
    Odrv4 I__6375 (
            .O(N__29871),
            .I(\QuadInstance0.Quad_RNO_0_0_2 ));
    InMux I__6374 (
            .O(N__29868),
            .I(\QuadInstance0.un1_Quad_cry_1 ));
    InMux I__6373 (
            .O(N__29865),
            .I(N__29862));
    LocalMux I__6372 (
            .O(N__29862),
            .I(N__29859));
    Span4Mux_h I__6371 (
            .O(N__29859),
            .I(N__29856));
    Span4Mux_h I__6370 (
            .O(N__29856),
            .I(N__29853));
    Odrv4 I__6369 (
            .O(N__29853),
            .I(\QuadInstance0.Quad_RNO_0_0_3 ));
    InMux I__6368 (
            .O(N__29850),
            .I(\QuadInstance0.un1_Quad_cry_2 ));
    InMux I__6367 (
            .O(N__29847),
            .I(N__29844));
    LocalMux I__6366 (
            .O(N__29844),
            .I(N__29841));
    Span4Mux_h I__6365 (
            .O(N__29841),
            .I(N__29838));
    Odrv4 I__6364 (
            .O(N__29838),
            .I(\QuadInstance0.Quad_RNO_0_0_4 ));
    InMux I__6363 (
            .O(N__29835),
            .I(\QuadInstance0.un1_Quad_cry_3 ));
    InMux I__6362 (
            .O(N__29832),
            .I(N__29829));
    LocalMux I__6361 (
            .O(N__29829),
            .I(N__29826));
    Odrv4 I__6360 (
            .O(N__29826),
            .I(\QuadInstance0.Quad_RNO_0_0_5 ));
    InMux I__6359 (
            .O(N__29823),
            .I(\QuadInstance0.un1_Quad_cry_4 ));
    InMux I__6358 (
            .O(N__29820),
            .I(N__29817));
    LocalMux I__6357 (
            .O(N__29817),
            .I(\PWMInstance3.un1_PWMPulseWidthCount_0_I_45_c_RNO_2 ));
    InMux I__6356 (
            .O(N__29814),
            .I(N__29811));
    LocalMux I__6355 (
            .O(N__29811),
            .I(N__29808));
    Odrv4 I__6354 (
            .O(N__29808),
            .I(\PWMInstance3.un1_PWMPulseWidthCount_0_I_33_c_RNO_2 ));
    InMux I__6353 (
            .O(N__29805),
            .I(N__29802));
    LocalMux I__6352 (
            .O(N__29802),
            .I(N__29799));
    Odrv4 I__6351 (
            .O(N__29799),
            .I(\PWMInstance3.un1_PWMPulseWidthCount_0_I_39_c_RNO_2 ));
    InMux I__6350 (
            .O(N__29796),
            .I(N__29793));
    LocalMux I__6349 (
            .O(N__29793),
            .I(N__29790));
    Odrv4 I__6348 (
            .O(N__29790),
            .I(\PWMInstance3.un1_PWMPulseWidthCount_0_I_21_c_RNO_2 ));
    InMux I__6347 (
            .O(N__29787),
            .I(N__29784));
    LocalMux I__6346 (
            .O(N__29784),
            .I(N__29781));
    Span4Mux_v I__6345 (
            .O(N__29781),
            .I(N__29778));
    Odrv4 I__6344 (
            .O(N__29778),
            .I(\PWMInstance3.un1_periodCounter12_1_0_a2_0 ));
    CascadeMux I__6343 (
            .O(N__29775),
            .I(N__29772));
    InMux I__6342 (
            .O(N__29772),
            .I(N__29768));
    InMux I__6341 (
            .O(N__29771),
            .I(N__29761));
    LocalMux I__6340 (
            .O(N__29768),
            .I(N__29758));
    InMux I__6339 (
            .O(N__29767),
            .I(N__29753));
    InMux I__6338 (
            .O(N__29766),
            .I(N__29753));
    InMux I__6337 (
            .O(N__29765),
            .I(N__29750));
    InMux I__6336 (
            .O(N__29764),
            .I(N__29747));
    LocalMux I__6335 (
            .O(N__29761),
            .I(N__29744));
    Span4Mux_h I__6334 (
            .O(N__29758),
            .I(N__29741));
    LocalMux I__6333 (
            .O(N__29753),
            .I(\PWMInstance3.out_0_sqmuxa ));
    LocalMux I__6332 (
            .O(N__29750),
            .I(\PWMInstance3.out_0_sqmuxa ));
    LocalMux I__6331 (
            .O(N__29747),
            .I(\PWMInstance3.out_0_sqmuxa ));
    Odrv4 I__6330 (
            .O(N__29744),
            .I(\PWMInstance3.out_0_sqmuxa ));
    Odrv4 I__6329 (
            .O(N__29741),
            .I(\PWMInstance3.out_0_sqmuxa ));
    InMux I__6328 (
            .O(N__29730),
            .I(bfn_16_16_0_));
    IoInMux I__6327 (
            .O(N__29727),
            .I(N__29724));
    LocalMux I__6326 (
            .O(N__29724),
            .I(N__29721));
    Span4Mux_s0_v I__6325 (
            .O(N__29721),
            .I(N__29718));
    Span4Mux_v I__6324 (
            .O(N__29718),
            .I(N__29714));
    InMux I__6323 (
            .O(N__29717),
            .I(N__29711));
    Odrv4 I__6322 (
            .O(N__29714),
            .I(PWM3_c));
    LocalMux I__6321 (
            .O(N__29711),
            .I(PWM3_c));
    InMux I__6320 (
            .O(N__29706),
            .I(N__29703));
    LocalMux I__6319 (
            .O(N__29703),
            .I(N__29700));
    IoSpan4Mux I__6318 (
            .O(N__29700),
            .I(N__29697));
    Odrv4 I__6317 (
            .O(N__29697),
            .I(ch7_A_c));
    InMux I__6316 (
            .O(N__29694),
            .I(N__29691));
    LocalMux I__6315 (
            .O(N__29691),
            .I(N__29688));
    Span4Mux_h I__6314 (
            .O(N__29688),
            .I(N__29685));
    Span4Mux_v I__6313 (
            .O(N__29685),
            .I(N__29682));
    Span4Mux_h I__6312 (
            .O(N__29682),
            .I(N__29679));
    Odrv4 I__6311 (
            .O(N__29679),
            .I(\QuadInstance7.delayedCh_AZ0Z_0 ));
    CascadeMux I__6310 (
            .O(N__29676),
            .I(N__29673));
    InMux I__6309 (
            .O(N__29673),
            .I(N__29670));
    LocalMux I__6308 (
            .O(N__29670),
            .I(N__29667));
    Odrv4 I__6307 (
            .O(N__29667),
            .I(\QuadInstance4.Quad_RNO_0_4_10 ));
    InMux I__6306 (
            .O(N__29664),
            .I(N__29653));
    InMux I__6305 (
            .O(N__29663),
            .I(N__29653));
    InMux I__6304 (
            .O(N__29662),
            .I(N__29649));
    InMux I__6303 (
            .O(N__29661),
            .I(N__29644));
    InMux I__6302 (
            .O(N__29660),
            .I(N__29644));
    InMux I__6301 (
            .O(N__29659),
            .I(N__29637));
    InMux I__6300 (
            .O(N__29658),
            .I(N__29637));
    LocalMux I__6299 (
            .O(N__29653),
            .I(N__29634));
    CascadeMux I__6298 (
            .O(N__29652),
            .I(N__29630));
    LocalMux I__6297 (
            .O(N__29649),
            .I(N__29625));
    LocalMux I__6296 (
            .O(N__29644),
            .I(N__29615));
    InMux I__6295 (
            .O(N__29643),
            .I(N__29610));
    InMux I__6294 (
            .O(N__29642),
            .I(N__29610));
    LocalMux I__6293 (
            .O(N__29637),
            .I(N__29605));
    Span4Mux_h I__6292 (
            .O(N__29634),
            .I(N__29605));
    InMux I__6291 (
            .O(N__29633),
            .I(N__29591));
    InMux I__6290 (
            .O(N__29630),
            .I(N__29591));
    InMux I__6289 (
            .O(N__29629),
            .I(N__29591));
    InMux I__6288 (
            .O(N__29628),
            .I(N__29584));
    Span4Mux_h I__6287 (
            .O(N__29625),
            .I(N__29581));
    InMux I__6286 (
            .O(N__29624),
            .I(N__29572));
    InMux I__6285 (
            .O(N__29623),
            .I(N__29572));
    InMux I__6284 (
            .O(N__29622),
            .I(N__29572));
    InMux I__6283 (
            .O(N__29621),
            .I(N__29572));
    InMux I__6282 (
            .O(N__29620),
            .I(N__29569));
    InMux I__6281 (
            .O(N__29619),
            .I(N__29564));
    InMux I__6280 (
            .O(N__29618),
            .I(N__29564));
    Span4Mux_v I__6279 (
            .O(N__29615),
            .I(N__29561));
    LocalMux I__6278 (
            .O(N__29610),
            .I(N__29556));
    Span4Mux_h I__6277 (
            .O(N__29605),
            .I(N__29556));
    InMux I__6276 (
            .O(N__29604),
            .I(N__29545));
    InMux I__6275 (
            .O(N__29603),
            .I(N__29545));
    InMux I__6274 (
            .O(N__29602),
            .I(N__29545));
    InMux I__6273 (
            .O(N__29601),
            .I(N__29545));
    InMux I__6272 (
            .O(N__29600),
            .I(N__29545));
    InMux I__6271 (
            .O(N__29599),
            .I(N__29540));
    InMux I__6270 (
            .O(N__29598),
            .I(N__29540));
    LocalMux I__6269 (
            .O(N__29591),
            .I(N__29537));
    InMux I__6268 (
            .O(N__29590),
            .I(N__29528));
    InMux I__6267 (
            .O(N__29589),
            .I(N__29528));
    InMux I__6266 (
            .O(N__29588),
            .I(N__29528));
    InMux I__6265 (
            .O(N__29587),
            .I(N__29528));
    LocalMux I__6264 (
            .O(N__29584),
            .I(N__29521));
    Span4Mux_h I__6263 (
            .O(N__29581),
            .I(N__29521));
    LocalMux I__6262 (
            .O(N__29572),
            .I(N__29521));
    LocalMux I__6261 (
            .O(N__29569),
            .I(quadWriteZ0Z_4));
    LocalMux I__6260 (
            .O(N__29564),
            .I(quadWriteZ0Z_4));
    Odrv4 I__6259 (
            .O(N__29561),
            .I(quadWriteZ0Z_4));
    Odrv4 I__6258 (
            .O(N__29556),
            .I(quadWriteZ0Z_4));
    LocalMux I__6257 (
            .O(N__29545),
            .I(quadWriteZ0Z_4));
    LocalMux I__6256 (
            .O(N__29540),
            .I(quadWriteZ0Z_4));
    Odrv4 I__6255 (
            .O(N__29537),
            .I(quadWriteZ0Z_4));
    LocalMux I__6254 (
            .O(N__29528),
            .I(quadWriteZ0Z_4));
    Odrv4 I__6253 (
            .O(N__29521),
            .I(quadWriteZ0Z_4));
    CascadeMux I__6252 (
            .O(N__29502),
            .I(N__29498));
    InMux I__6251 (
            .O(N__29501),
            .I(N__29494));
    InMux I__6250 (
            .O(N__29498),
            .I(N__29491));
    InMux I__6249 (
            .O(N__29497),
            .I(N__29488));
    LocalMux I__6248 (
            .O(N__29494),
            .I(\PWMInstance3.periodCounterZ0Z_7 ));
    LocalMux I__6247 (
            .O(N__29491),
            .I(\PWMInstance3.periodCounterZ0Z_7 ));
    LocalMux I__6246 (
            .O(N__29488),
            .I(\PWMInstance3.periodCounterZ0Z_7 ));
    InMux I__6245 (
            .O(N__29481),
            .I(N__29476));
    InMux I__6244 (
            .O(N__29480),
            .I(N__29471));
    InMux I__6243 (
            .O(N__29479),
            .I(N__29471));
    LocalMux I__6242 (
            .O(N__29476),
            .I(\PWMInstance3.periodCounterZ0Z_6 ));
    LocalMux I__6241 (
            .O(N__29471),
            .I(\PWMInstance3.periodCounterZ0Z_6 ));
    InMux I__6240 (
            .O(N__29466),
            .I(N__29463));
    LocalMux I__6239 (
            .O(N__29463),
            .I(\PWMInstance3.PWMPulseWidthCountZ0Z_6 ));
    InMux I__6238 (
            .O(N__29460),
            .I(N__29457));
    LocalMux I__6237 (
            .O(N__29457),
            .I(N__29453));
    InMux I__6236 (
            .O(N__29456),
            .I(N__29445));
    Span4Mux_v I__6235 (
            .O(N__29453),
            .I(N__29440));
    InMux I__6234 (
            .O(N__29452),
            .I(N__29431));
    InMux I__6233 (
            .O(N__29451),
            .I(N__29431));
    InMux I__6232 (
            .O(N__29450),
            .I(N__29431));
    InMux I__6231 (
            .O(N__29449),
            .I(N__29431));
    InMux I__6230 (
            .O(N__29448),
            .I(N__29428));
    LocalMux I__6229 (
            .O(N__29445),
            .I(N__29422));
    InMux I__6228 (
            .O(N__29444),
            .I(N__29419));
    CascadeMux I__6227 (
            .O(N__29443),
            .I(N__29414));
    Span4Mux_h I__6226 (
            .O(N__29440),
            .I(N__29406));
    LocalMux I__6225 (
            .O(N__29431),
            .I(N__29406));
    LocalMux I__6224 (
            .O(N__29428),
            .I(N__29406));
    InMux I__6223 (
            .O(N__29427),
            .I(N__29401));
    InMux I__6222 (
            .O(N__29426),
            .I(N__29401));
    InMux I__6221 (
            .O(N__29425),
            .I(N__29398));
    Span4Mux_h I__6220 (
            .O(N__29422),
            .I(N__29393));
    LocalMux I__6219 (
            .O(N__29419),
            .I(N__29393));
    InMux I__6218 (
            .O(N__29418),
            .I(N__29389));
    InMux I__6217 (
            .O(N__29417),
            .I(N__29386));
    InMux I__6216 (
            .O(N__29414),
            .I(N__29383));
    InMux I__6215 (
            .O(N__29413),
            .I(N__29380));
    Span4Mux_h I__6214 (
            .O(N__29406),
            .I(N__29375));
    LocalMux I__6213 (
            .O(N__29401),
            .I(N__29375));
    LocalMux I__6212 (
            .O(N__29398),
            .I(N__29372));
    Span4Mux_h I__6211 (
            .O(N__29393),
            .I(N__29369));
    InMux I__6210 (
            .O(N__29392),
            .I(N__29366));
    LocalMux I__6209 (
            .O(N__29389),
            .I(N__29363));
    LocalMux I__6208 (
            .O(N__29386),
            .I(N__29358));
    LocalMux I__6207 (
            .O(N__29383),
            .I(N__29358));
    LocalMux I__6206 (
            .O(N__29380),
            .I(N__29355));
    Span4Mux_h I__6205 (
            .O(N__29375),
            .I(N__29352));
    Span4Mux_h I__6204 (
            .O(N__29372),
            .I(N__29349));
    Span4Mux_v I__6203 (
            .O(N__29369),
            .I(N__29344));
    LocalMux I__6202 (
            .O(N__29366),
            .I(N__29344));
    Span12Mux_s11_h I__6201 (
            .O(N__29363),
            .I(N__29339));
    Span12Mux_h I__6200 (
            .O(N__29358),
            .I(N__29339));
    Span4Mux_h I__6199 (
            .O(N__29355),
            .I(N__29334));
    Span4Mux_v I__6198 (
            .O(N__29352),
            .I(N__29334));
    Odrv4 I__6197 (
            .O(N__29349),
            .I(dataWriteZ0Z_7));
    Odrv4 I__6196 (
            .O(N__29344),
            .I(dataWriteZ0Z_7));
    Odrv12 I__6195 (
            .O(N__29339),
            .I(dataWriteZ0Z_7));
    Odrv4 I__6194 (
            .O(N__29334),
            .I(dataWriteZ0Z_7));
    InMux I__6193 (
            .O(N__29325),
            .I(N__29322));
    LocalMux I__6192 (
            .O(N__29322),
            .I(\PWMInstance3.PWMPulseWidthCountZ0Z_7 ));
    CEMux I__6191 (
            .O(N__29319),
            .I(N__29315));
    CEMux I__6190 (
            .O(N__29318),
            .I(N__29312));
    LocalMux I__6189 (
            .O(N__29315),
            .I(N__29309));
    LocalMux I__6188 (
            .O(N__29312),
            .I(N__29305));
    Span4Mux_v I__6187 (
            .O(N__29309),
            .I(N__29302));
    CEMux I__6186 (
            .O(N__29308),
            .I(N__29299));
    Span4Mux_v I__6185 (
            .O(N__29305),
            .I(N__29291));
    Span4Mux_v I__6184 (
            .O(N__29302),
            .I(N__29291));
    LocalMux I__6183 (
            .O(N__29299),
            .I(N__29291));
    CEMux I__6182 (
            .O(N__29298),
            .I(N__29287));
    Span4Mux_v I__6181 (
            .O(N__29291),
            .I(N__29284));
    CEMux I__6180 (
            .O(N__29290),
            .I(N__29281));
    LocalMux I__6179 (
            .O(N__29287),
            .I(\PWMInstance3.pwmWrite_0_3 ));
    Odrv4 I__6178 (
            .O(N__29284),
            .I(\PWMInstance3.pwmWrite_0_3 ));
    LocalMux I__6177 (
            .O(N__29281),
            .I(\PWMInstance3.pwmWrite_0_3 ));
    InMux I__6176 (
            .O(N__29274),
            .I(N__29271));
    LocalMux I__6175 (
            .O(N__29271),
            .I(N__29268));
    Span4Mux_v I__6174 (
            .O(N__29268),
            .I(N__29265));
    Odrv4 I__6173 (
            .O(N__29265),
            .I(\PWMInstance3.PWMPulseWidthCountZ0Z_8 ));
    CascadeMux I__6172 (
            .O(N__29262),
            .I(N__29258));
    InMux I__6171 (
            .O(N__29261),
            .I(N__29254));
    InMux I__6170 (
            .O(N__29258),
            .I(N__29249));
    InMux I__6169 (
            .O(N__29257),
            .I(N__29249));
    LocalMux I__6168 (
            .O(N__29254),
            .I(\PWMInstance3.periodCounterZ0Z_8 ));
    LocalMux I__6167 (
            .O(N__29249),
            .I(\PWMInstance3.periodCounterZ0Z_8 ));
    CascadeMux I__6166 (
            .O(N__29244),
            .I(N__29239));
    InMux I__6165 (
            .O(N__29243),
            .I(N__29236));
    InMux I__6164 (
            .O(N__29242),
            .I(N__29233));
    InMux I__6163 (
            .O(N__29239),
            .I(N__29230));
    LocalMux I__6162 (
            .O(N__29236),
            .I(\PWMInstance3.periodCounterZ0Z_9 ));
    LocalMux I__6161 (
            .O(N__29233),
            .I(\PWMInstance3.periodCounterZ0Z_9 ));
    LocalMux I__6160 (
            .O(N__29230),
            .I(\PWMInstance3.periodCounterZ0Z_9 ));
    InMux I__6159 (
            .O(N__29223),
            .I(N__29220));
    LocalMux I__6158 (
            .O(N__29220),
            .I(N__29217));
    Odrv4 I__6157 (
            .O(N__29217),
            .I(\PWMInstance3.PWMPulseWidthCountZ0Z_9 ));
    InMux I__6156 (
            .O(N__29214),
            .I(N__29211));
    LocalMux I__6155 (
            .O(N__29211),
            .I(\PWMInstance3.un1_PWMPulseWidthCount_0_I_1_c_RNO_2 ));
    InMux I__6154 (
            .O(N__29208),
            .I(N__29205));
    LocalMux I__6153 (
            .O(N__29205),
            .I(N__29202));
    Odrv4 I__6152 (
            .O(N__29202),
            .I(\PWMInstance3.un1_PWMPulseWidthCount_0_I_9_c_RNO_2 ));
    InMux I__6151 (
            .O(N__29199),
            .I(N__29196));
    LocalMux I__6150 (
            .O(N__29196),
            .I(N__29193));
    Span4Mux_v I__6149 (
            .O(N__29193),
            .I(N__29190));
    Odrv4 I__6148 (
            .O(N__29190),
            .I(\PWMInstance3.un1_PWMPulseWidthCount_0_I_15_c_RNO_2 ));
    InMux I__6147 (
            .O(N__29187),
            .I(N__29184));
    LocalMux I__6146 (
            .O(N__29184),
            .I(\PWMInstance3.un1_PWMPulseWidthCount_0_I_27_c_RNO_2 ));
    InMux I__6145 (
            .O(N__29181),
            .I(N__29178));
    LocalMux I__6144 (
            .O(N__29178),
            .I(\PWMInstance3.PWMPulseWidthCountZ0Z_2 ));
    CascadeMux I__6143 (
            .O(N__29175),
            .I(N__29171));
    InMux I__6142 (
            .O(N__29174),
            .I(N__29167));
    InMux I__6141 (
            .O(N__29171),
            .I(N__29164));
    InMux I__6140 (
            .O(N__29170),
            .I(N__29161));
    LocalMux I__6139 (
            .O(N__29167),
            .I(\PWMInstance3.periodCounterZ0Z_15 ));
    LocalMux I__6138 (
            .O(N__29164),
            .I(\PWMInstance3.periodCounterZ0Z_15 ));
    LocalMux I__6137 (
            .O(N__29161),
            .I(\PWMInstance3.periodCounterZ0Z_15 ));
    InMux I__6136 (
            .O(N__29154),
            .I(N__29149));
    InMux I__6135 (
            .O(N__29153),
            .I(N__29146));
    InMux I__6134 (
            .O(N__29152),
            .I(N__29143));
    LocalMux I__6133 (
            .O(N__29149),
            .I(N__29140));
    LocalMux I__6132 (
            .O(N__29146),
            .I(\PWMInstance3.periodCounterZ0Z_14 ));
    LocalMux I__6131 (
            .O(N__29143),
            .I(\PWMInstance3.periodCounterZ0Z_14 ));
    Odrv4 I__6130 (
            .O(N__29140),
            .I(\PWMInstance3.periodCounterZ0Z_14 ));
    InMux I__6129 (
            .O(N__29133),
            .I(N__29130));
    LocalMux I__6128 (
            .O(N__29130),
            .I(\PWMInstance3.PWMPulseWidthCountZ0Z_14 ));
    InMux I__6127 (
            .O(N__29127),
            .I(N__29124));
    LocalMux I__6126 (
            .O(N__29124),
            .I(\PWMInstance3.PWMPulseWidthCountZ0Z_15 ));
    InMux I__6125 (
            .O(N__29121),
            .I(N__29118));
    LocalMux I__6124 (
            .O(N__29118),
            .I(\PWMInstance3.PWMPulseWidthCountZ0Z_13 ));
    InMux I__6123 (
            .O(N__29115),
            .I(N__29112));
    LocalMux I__6122 (
            .O(N__29112),
            .I(\PWMInstance3.PWMPulseWidthCountZ0Z_12 ));
    InMux I__6121 (
            .O(N__29109),
            .I(N__29104));
    InMux I__6120 (
            .O(N__29108),
            .I(N__29101));
    InMux I__6119 (
            .O(N__29107),
            .I(N__29098));
    LocalMux I__6118 (
            .O(N__29104),
            .I(N__29095));
    LocalMux I__6117 (
            .O(N__29101),
            .I(\PWMInstance3.periodCounterZ0Z_12 ));
    LocalMux I__6116 (
            .O(N__29098),
            .I(\PWMInstance3.periodCounterZ0Z_12 ));
    Odrv4 I__6115 (
            .O(N__29095),
            .I(\PWMInstance3.periodCounterZ0Z_12 ));
    CascadeMux I__6114 (
            .O(N__29088),
            .I(N__29084));
    InMux I__6113 (
            .O(N__29087),
            .I(N__29080));
    InMux I__6112 (
            .O(N__29084),
            .I(N__29077));
    InMux I__6111 (
            .O(N__29083),
            .I(N__29074));
    LocalMux I__6110 (
            .O(N__29080),
            .I(\PWMInstance3.periodCounterZ0Z_13 ));
    LocalMux I__6109 (
            .O(N__29077),
            .I(\PWMInstance3.periodCounterZ0Z_13 ));
    LocalMux I__6108 (
            .O(N__29074),
            .I(\PWMInstance3.periodCounterZ0Z_13 ));
    InMux I__6107 (
            .O(N__29067),
            .I(N__29064));
    LocalMux I__6106 (
            .O(N__29064),
            .I(N__29061));
    Span4Mux_v I__6105 (
            .O(N__29061),
            .I(N__29058));
    Odrv4 I__6104 (
            .O(N__29058),
            .I(\PWMInstance3.un1_periodCounter12_1_0_a2_0_9 ));
    InMux I__6103 (
            .O(N__29055),
            .I(N__29050));
    InMux I__6102 (
            .O(N__29054),
            .I(N__29045));
    InMux I__6101 (
            .O(N__29053),
            .I(N__29045));
    LocalMux I__6100 (
            .O(N__29050),
            .I(\PWMInstance3.periodCounterZ0Z_0 ));
    LocalMux I__6099 (
            .O(N__29045),
            .I(\PWMInstance3.periodCounterZ0Z_0 ));
    CascadeMux I__6098 (
            .O(N__29040),
            .I(N__29035));
    InMux I__6097 (
            .O(N__29039),
            .I(N__29032));
    InMux I__6096 (
            .O(N__29038),
            .I(N__29029));
    InMux I__6095 (
            .O(N__29035),
            .I(N__29026));
    LocalMux I__6094 (
            .O(N__29032),
            .I(\PWMInstance3.periodCounterZ0Z_1 ));
    LocalMux I__6093 (
            .O(N__29029),
            .I(\PWMInstance3.periodCounterZ0Z_1 ));
    LocalMux I__6092 (
            .O(N__29026),
            .I(\PWMInstance3.periodCounterZ0Z_1 ));
    InMux I__6091 (
            .O(N__29019),
            .I(N__29016));
    LocalMux I__6090 (
            .O(N__29016),
            .I(\PWMInstance3.PWMPulseWidthCountZ0Z_0 ));
    InMux I__6089 (
            .O(N__29013),
            .I(N__29010));
    LocalMux I__6088 (
            .O(N__29010),
            .I(\PWMInstance3.PWMPulseWidthCountZ0Z_1 ));
    InMux I__6087 (
            .O(N__29007),
            .I(N__29004));
    LocalMux I__6086 (
            .O(N__29004),
            .I(N__28999));
    InMux I__6085 (
            .O(N__29003),
            .I(N__28996));
    InMux I__6084 (
            .O(N__29002),
            .I(N__28993));
    Span4Mux_v I__6083 (
            .O(N__28999),
            .I(N__28980));
    LocalMux I__6082 (
            .O(N__28996),
            .I(N__28980));
    LocalMux I__6081 (
            .O(N__28993),
            .I(N__28977));
    InMux I__6080 (
            .O(N__28992),
            .I(N__28973));
    InMux I__6079 (
            .O(N__28991),
            .I(N__28967));
    InMux I__6078 (
            .O(N__28990),
            .I(N__28967));
    InMux I__6077 (
            .O(N__28989),
            .I(N__28962));
    InMux I__6076 (
            .O(N__28988),
            .I(N__28962));
    InMux I__6075 (
            .O(N__28987),
            .I(N__28959));
    InMux I__6074 (
            .O(N__28986),
            .I(N__28956));
    InMux I__6073 (
            .O(N__28985),
            .I(N__28953));
    Span4Mux_v I__6072 (
            .O(N__28980),
            .I(N__28947));
    Span4Mux_v I__6071 (
            .O(N__28977),
            .I(N__28947));
    InMux I__6070 (
            .O(N__28976),
            .I(N__28944));
    LocalMux I__6069 (
            .O(N__28973),
            .I(N__28940));
    InMux I__6068 (
            .O(N__28972),
            .I(N__28937));
    LocalMux I__6067 (
            .O(N__28967),
            .I(N__28934));
    LocalMux I__6066 (
            .O(N__28962),
            .I(N__28925));
    LocalMux I__6065 (
            .O(N__28959),
            .I(N__28925));
    LocalMux I__6064 (
            .O(N__28956),
            .I(N__28925));
    LocalMux I__6063 (
            .O(N__28953),
            .I(N__28925));
    InMux I__6062 (
            .O(N__28952),
            .I(N__28922));
    Span4Mux_h I__6061 (
            .O(N__28947),
            .I(N__28919));
    LocalMux I__6060 (
            .O(N__28944),
            .I(N__28916));
    InMux I__6059 (
            .O(N__28943),
            .I(N__28913));
    Span4Mux_v I__6058 (
            .O(N__28940),
            .I(N__28909));
    LocalMux I__6057 (
            .O(N__28937),
            .I(N__28904));
    Span4Mux_v I__6056 (
            .O(N__28934),
            .I(N__28904));
    Span4Mux_v I__6055 (
            .O(N__28925),
            .I(N__28899));
    LocalMux I__6054 (
            .O(N__28922),
            .I(N__28899));
    Span4Mux_h I__6053 (
            .O(N__28919),
            .I(N__28892));
    Span4Mux_v I__6052 (
            .O(N__28916),
            .I(N__28892));
    LocalMux I__6051 (
            .O(N__28913),
            .I(N__28892));
    InMux I__6050 (
            .O(N__28912),
            .I(N__28889));
    Span4Mux_h I__6049 (
            .O(N__28909),
            .I(N__28882));
    Span4Mux_v I__6048 (
            .O(N__28904),
            .I(N__28882));
    Span4Mux_v I__6047 (
            .O(N__28899),
            .I(N__28882));
    Odrv4 I__6046 (
            .O(N__28892),
            .I(dataWriteZ0Z_8));
    LocalMux I__6045 (
            .O(N__28889),
            .I(dataWriteZ0Z_8));
    Odrv4 I__6044 (
            .O(N__28882),
            .I(dataWriteZ0Z_8));
    InMux I__6043 (
            .O(N__28875),
            .I(N__28867));
    CascadeMux I__6042 (
            .O(N__28874),
            .I(N__28863));
    InMux I__6041 (
            .O(N__28873),
            .I(N__28858));
    InMux I__6040 (
            .O(N__28872),
            .I(N__28855));
    InMux I__6039 (
            .O(N__28871),
            .I(N__28851));
    InMux I__6038 (
            .O(N__28870),
            .I(N__28848));
    LocalMux I__6037 (
            .O(N__28867),
            .I(N__28844));
    InMux I__6036 (
            .O(N__28866),
            .I(N__28839));
    InMux I__6035 (
            .O(N__28863),
            .I(N__28839));
    InMux I__6034 (
            .O(N__28862),
            .I(N__28834));
    InMux I__6033 (
            .O(N__28861),
            .I(N__28834));
    LocalMux I__6032 (
            .O(N__28858),
            .I(N__28830));
    LocalMux I__6031 (
            .O(N__28855),
            .I(N__28827));
    InMux I__6030 (
            .O(N__28854),
            .I(N__28824));
    LocalMux I__6029 (
            .O(N__28851),
            .I(N__28820));
    LocalMux I__6028 (
            .O(N__28848),
            .I(N__28816));
    InMux I__6027 (
            .O(N__28847),
            .I(N__28813));
    Span4Mux_v I__6026 (
            .O(N__28844),
            .I(N__28808));
    LocalMux I__6025 (
            .O(N__28839),
            .I(N__28808));
    LocalMux I__6024 (
            .O(N__28834),
            .I(N__28805));
    InMux I__6023 (
            .O(N__28833),
            .I(N__28802));
    Span4Mux_h I__6022 (
            .O(N__28830),
            .I(N__28797));
    Span4Mux_h I__6021 (
            .O(N__28827),
            .I(N__28794));
    LocalMux I__6020 (
            .O(N__28824),
            .I(N__28791));
    InMux I__6019 (
            .O(N__28823),
            .I(N__28788));
    Span4Mux_v I__6018 (
            .O(N__28820),
            .I(N__28785));
    InMux I__6017 (
            .O(N__28819),
            .I(N__28782));
    Span4Mux_v I__6016 (
            .O(N__28816),
            .I(N__28779));
    LocalMux I__6015 (
            .O(N__28813),
            .I(N__28776));
    Span4Mux_h I__6014 (
            .O(N__28808),
            .I(N__28769));
    Span4Mux_h I__6013 (
            .O(N__28805),
            .I(N__28769));
    LocalMux I__6012 (
            .O(N__28802),
            .I(N__28769));
    InMux I__6011 (
            .O(N__28801),
            .I(N__28766));
    InMux I__6010 (
            .O(N__28800),
            .I(N__28763));
    Span4Mux_h I__6009 (
            .O(N__28797),
            .I(N__28760));
    Span4Mux_h I__6008 (
            .O(N__28794),
            .I(N__28753));
    Span4Mux_v I__6007 (
            .O(N__28791),
            .I(N__28753));
    LocalMux I__6006 (
            .O(N__28788),
            .I(N__28753));
    Sp12to4 I__6005 (
            .O(N__28785),
            .I(N__28748));
    LocalMux I__6004 (
            .O(N__28782),
            .I(N__28748));
    Span4Mux_h I__6003 (
            .O(N__28779),
            .I(N__28737));
    Span4Mux_h I__6002 (
            .O(N__28776),
            .I(N__28737));
    Span4Mux_h I__6001 (
            .O(N__28769),
            .I(N__28737));
    LocalMux I__6000 (
            .O(N__28766),
            .I(N__28737));
    LocalMux I__5999 (
            .O(N__28763),
            .I(N__28737));
    Odrv4 I__5998 (
            .O(N__28760),
            .I(dataWriteZ0Z_12));
    Odrv4 I__5997 (
            .O(N__28753),
            .I(dataWriteZ0Z_12));
    Odrv12 I__5996 (
            .O(N__28748),
            .I(dataWriteZ0Z_12));
    Odrv4 I__5995 (
            .O(N__28737),
            .I(dataWriteZ0Z_12));
    InMux I__5994 (
            .O(N__28728),
            .I(N__28720));
    InMux I__5993 (
            .O(N__28727),
            .I(N__28716));
    InMux I__5992 (
            .O(N__28726),
            .I(N__28712));
    InMux I__5991 (
            .O(N__28725),
            .I(N__28708));
    InMux I__5990 (
            .O(N__28724),
            .I(N__28705));
    InMux I__5989 (
            .O(N__28723),
            .I(N__28700));
    LocalMux I__5988 (
            .O(N__28720),
            .I(N__28696));
    InMux I__5987 (
            .O(N__28719),
            .I(N__28693));
    LocalMux I__5986 (
            .O(N__28716),
            .I(N__28690));
    InMux I__5985 (
            .O(N__28715),
            .I(N__28687));
    LocalMux I__5984 (
            .O(N__28712),
            .I(N__28681));
    InMux I__5983 (
            .O(N__28711),
            .I(N__28678));
    LocalMux I__5982 (
            .O(N__28708),
            .I(N__28674));
    LocalMux I__5981 (
            .O(N__28705),
            .I(N__28671));
    InMux I__5980 (
            .O(N__28704),
            .I(N__28668));
    InMux I__5979 (
            .O(N__28703),
            .I(N__28665));
    LocalMux I__5978 (
            .O(N__28700),
            .I(N__28662));
    InMux I__5977 (
            .O(N__28699),
            .I(N__28659));
    Span4Mux_v I__5976 (
            .O(N__28696),
            .I(N__28654));
    LocalMux I__5975 (
            .O(N__28693),
            .I(N__28654));
    Span4Mux_h I__5974 (
            .O(N__28690),
            .I(N__28649));
    LocalMux I__5973 (
            .O(N__28687),
            .I(N__28649));
    InMux I__5972 (
            .O(N__28686),
            .I(N__28642));
    InMux I__5971 (
            .O(N__28685),
            .I(N__28642));
    InMux I__5970 (
            .O(N__28684),
            .I(N__28642));
    Span4Mux_v I__5969 (
            .O(N__28681),
            .I(N__28639));
    LocalMux I__5968 (
            .O(N__28678),
            .I(N__28636));
    InMux I__5967 (
            .O(N__28677),
            .I(N__28633));
    Span4Mux_h I__5966 (
            .O(N__28674),
            .I(N__28630));
    Span4Mux_v I__5965 (
            .O(N__28671),
            .I(N__28623));
    LocalMux I__5964 (
            .O(N__28668),
            .I(N__28623));
    LocalMux I__5963 (
            .O(N__28665),
            .I(N__28623));
    Span4Mux_v I__5962 (
            .O(N__28662),
            .I(N__28620));
    LocalMux I__5961 (
            .O(N__28659),
            .I(N__28617));
    Span4Mux_h I__5960 (
            .O(N__28654),
            .I(N__28610));
    Span4Mux_h I__5959 (
            .O(N__28649),
            .I(N__28610));
    LocalMux I__5958 (
            .O(N__28642),
            .I(N__28610));
    Span4Mux_h I__5957 (
            .O(N__28639),
            .I(N__28603));
    Span4Mux_v I__5956 (
            .O(N__28636),
            .I(N__28603));
    LocalMux I__5955 (
            .O(N__28633),
            .I(N__28603));
    Span4Mux_h I__5954 (
            .O(N__28630),
            .I(N__28598));
    Span4Mux_h I__5953 (
            .O(N__28623),
            .I(N__28598));
    Span4Mux_h I__5952 (
            .O(N__28620),
            .I(N__28591));
    Span4Mux_h I__5951 (
            .O(N__28617),
            .I(N__28591));
    Span4Mux_v I__5950 (
            .O(N__28610),
            .I(N__28591));
    Odrv4 I__5949 (
            .O(N__28603),
            .I(dataWriteZ0Z_13));
    Odrv4 I__5948 (
            .O(N__28598),
            .I(dataWriteZ0Z_13));
    Odrv4 I__5947 (
            .O(N__28591),
            .I(dataWriteZ0Z_13));
    InMux I__5946 (
            .O(N__28584),
            .I(N__28581));
    LocalMux I__5945 (
            .O(N__28581),
            .I(N__28573));
    InMux I__5944 (
            .O(N__28580),
            .I(N__28569));
    InMux I__5943 (
            .O(N__28579),
            .I(N__28566));
    InMux I__5942 (
            .O(N__28578),
            .I(N__28560));
    InMux I__5941 (
            .O(N__28577),
            .I(N__28560));
    InMux I__5940 (
            .O(N__28576),
            .I(N__28554));
    Span4Mux_v I__5939 (
            .O(N__28573),
            .I(N__28551));
    InMux I__5938 (
            .O(N__28572),
            .I(N__28548));
    LocalMux I__5937 (
            .O(N__28569),
            .I(N__28545));
    LocalMux I__5936 (
            .O(N__28566),
            .I(N__28542));
    InMux I__5935 (
            .O(N__28565),
            .I(N__28538));
    LocalMux I__5934 (
            .O(N__28560),
            .I(N__28535));
    InMux I__5933 (
            .O(N__28559),
            .I(N__28532));
    InMux I__5932 (
            .O(N__28558),
            .I(N__28529));
    InMux I__5931 (
            .O(N__28557),
            .I(N__28524));
    LocalMux I__5930 (
            .O(N__28554),
            .I(N__28520));
    Span4Mux_h I__5929 (
            .O(N__28551),
            .I(N__28515));
    LocalMux I__5928 (
            .O(N__28548),
            .I(N__28515));
    Span4Mux_v I__5927 (
            .O(N__28545),
            .I(N__28510));
    Span4Mux_v I__5926 (
            .O(N__28542),
            .I(N__28510));
    InMux I__5925 (
            .O(N__28541),
            .I(N__28507));
    LocalMux I__5924 (
            .O(N__28538),
            .I(N__28503));
    Span4Mux_h I__5923 (
            .O(N__28535),
            .I(N__28496));
    LocalMux I__5922 (
            .O(N__28532),
            .I(N__28496));
    LocalMux I__5921 (
            .O(N__28529),
            .I(N__28496));
    InMux I__5920 (
            .O(N__28528),
            .I(N__28491));
    InMux I__5919 (
            .O(N__28527),
            .I(N__28491));
    LocalMux I__5918 (
            .O(N__28524),
            .I(N__28488));
    InMux I__5917 (
            .O(N__28523),
            .I(N__28485));
    Span4Mux_h I__5916 (
            .O(N__28520),
            .I(N__28482));
    Span4Mux_h I__5915 (
            .O(N__28515),
            .I(N__28479));
    Span4Mux_h I__5914 (
            .O(N__28510),
            .I(N__28476));
    LocalMux I__5913 (
            .O(N__28507),
            .I(N__28473));
    InMux I__5912 (
            .O(N__28506),
            .I(N__28470));
    Span4Mux_v I__5911 (
            .O(N__28503),
            .I(N__28463));
    Span4Mux_h I__5910 (
            .O(N__28496),
            .I(N__28463));
    LocalMux I__5909 (
            .O(N__28491),
            .I(N__28463));
    Span4Mux_v I__5908 (
            .O(N__28488),
            .I(N__28458));
    LocalMux I__5907 (
            .O(N__28485),
            .I(N__28458));
    Span4Mux_h I__5906 (
            .O(N__28482),
            .I(N__28453));
    Span4Mux_v I__5905 (
            .O(N__28479),
            .I(N__28453));
    Span4Mux_h I__5904 (
            .O(N__28476),
            .I(N__28444));
    Span4Mux_v I__5903 (
            .O(N__28473),
            .I(N__28444));
    LocalMux I__5902 (
            .O(N__28470),
            .I(N__28444));
    Span4Mux_v I__5901 (
            .O(N__28463),
            .I(N__28444));
    Odrv4 I__5900 (
            .O(N__28458),
            .I(dataWriteZ0Z_9));
    Odrv4 I__5899 (
            .O(N__28453),
            .I(dataWriteZ0Z_9));
    Odrv4 I__5898 (
            .O(N__28444),
            .I(dataWriteZ0Z_9));
    CascadeMux I__5897 (
            .O(N__28437),
            .I(N__28432));
    InMux I__5896 (
            .O(N__28436),
            .I(N__28429));
    InMux I__5895 (
            .O(N__28435),
            .I(N__28426));
    InMux I__5894 (
            .O(N__28432),
            .I(N__28423));
    LocalMux I__5893 (
            .O(N__28429),
            .I(\PWMInstance3.periodCounterZ0Z_5 ));
    LocalMux I__5892 (
            .O(N__28426),
            .I(\PWMInstance3.periodCounterZ0Z_5 ));
    LocalMux I__5891 (
            .O(N__28423),
            .I(\PWMInstance3.periodCounterZ0Z_5 ));
    CascadeMux I__5890 (
            .O(N__28416),
            .I(N__28412));
    CascadeMux I__5889 (
            .O(N__28415),
            .I(N__28408));
    InMux I__5888 (
            .O(N__28412),
            .I(N__28405));
    InMux I__5887 (
            .O(N__28411),
            .I(N__28402));
    InMux I__5886 (
            .O(N__28408),
            .I(N__28399));
    LocalMux I__5885 (
            .O(N__28405),
            .I(N__28396));
    LocalMux I__5884 (
            .O(N__28402),
            .I(\PWMInstance3.periodCounterZ0Z_11 ));
    LocalMux I__5883 (
            .O(N__28399),
            .I(\PWMInstance3.periodCounterZ0Z_11 ));
    Odrv4 I__5882 (
            .O(N__28396),
            .I(\PWMInstance3.periodCounterZ0Z_11 ));
    InMux I__5881 (
            .O(N__28389),
            .I(N__28386));
    LocalMux I__5880 (
            .O(N__28386),
            .I(N__28383));
    Odrv4 I__5879 (
            .O(N__28383),
            .I(\PWMInstance3.un1_periodCounter12_1_0_a2_0_10 ));
    InMux I__5878 (
            .O(N__28380),
            .I(N__28377));
    LocalMux I__5877 (
            .O(N__28377),
            .I(N__28374));
    Span4Mux_h I__5876 (
            .O(N__28374),
            .I(N__28371));
    Odrv4 I__5875 (
            .O(N__28371),
            .I(\PWMInstance3.PWMPulseWidthCountZ0Z_3 ));
    CascadeMux I__5874 (
            .O(N__28368),
            .I(N__28363));
    InMux I__5873 (
            .O(N__28367),
            .I(N__28360));
    InMux I__5872 (
            .O(N__28366),
            .I(N__28355));
    InMux I__5871 (
            .O(N__28363),
            .I(N__28355));
    LocalMux I__5870 (
            .O(N__28360),
            .I(\PWMInstance3.periodCounterZ0Z_3 ));
    LocalMux I__5869 (
            .O(N__28355),
            .I(\PWMInstance3.periodCounterZ0Z_3 ));
    InMux I__5868 (
            .O(N__28350),
            .I(N__28345));
    InMux I__5867 (
            .O(N__28349),
            .I(N__28342));
    InMux I__5866 (
            .O(N__28348),
            .I(N__28339));
    LocalMux I__5865 (
            .O(N__28345),
            .I(\PWMInstance3.periodCounterZ0Z_2 ));
    LocalMux I__5864 (
            .O(N__28342),
            .I(\PWMInstance3.periodCounterZ0Z_2 ));
    LocalMux I__5863 (
            .O(N__28339),
            .I(\PWMInstance3.periodCounterZ0Z_2 ));
    CascadeMux I__5862 (
            .O(N__28332),
            .I(OutReg_esr_RNO_1Z0Z_6_cascade_));
    InMux I__5861 (
            .O(N__28329),
            .I(N__28326));
    LocalMux I__5860 (
            .O(N__28326),
            .I(N__28323));
    Span4Mux_v I__5859 (
            .O(N__28323),
            .I(N__28320));
    Odrv4 I__5858 (
            .O(N__28320),
            .I(OutReg_esr_RNO_2Z0Z_6));
    CascadeMux I__5857 (
            .O(N__28317),
            .I(OutReg_esr_RNO_0Z0Z_6_cascade_));
    InMux I__5856 (
            .O(N__28314),
            .I(N__28311));
    LocalMux I__5855 (
            .O(N__28311),
            .I(N__28308));
    Odrv4 I__5854 (
            .O(N__28308),
            .I(OutRegZ0Z_6));
    InMux I__5853 (
            .O(N__28305),
            .I(N__28301));
    InMux I__5852 (
            .O(N__28304),
            .I(N__28297));
    LocalMux I__5851 (
            .O(N__28301),
            .I(N__28294));
    InMux I__5850 (
            .O(N__28300),
            .I(N__28291));
    LocalMux I__5849 (
            .O(N__28297),
            .I(N__28288));
    Span4Mux_v I__5848 (
            .O(N__28294),
            .I(N__28283));
    LocalMux I__5847 (
            .O(N__28291),
            .I(N__28283));
    Span4Mux_v I__5846 (
            .O(N__28288),
            .I(N__28280));
    Span4Mux_v I__5845 (
            .O(N__28283),
            .I(N__28277));
    Span4Mux_h I__5844 (
            .O(N__28280),
            .I(N__28274));
    Odrv4 I__5843 (
            .O(N__28277),
            .I(dataRead2_6));
    Odrv4 I__5842 (
            .O(N__28274),
            .I(dataRead2_6));
    CascadeMux I__5841 (
            .O(N__28269),
            .I(N__28266));
    InMux I__5840 (
            .O(N__28266),
            .I(N__28262));
    InMux I__5839 (
            .O(N__28265),
            .I(N__28259));
    LocalMux I__5838 (
            .O(N__28262),
            .I(N__28255));
    LocalMux I__5837 (
            .O(N__28259),
            .I(N__28252));
    InMux I__5836 (
            .O(N__28258),
            .I(N__28249));
    Span4Mux_v I__5835 (
            .O(N__28255),
            .I(N__28246));
    Span4Mux_v I__5834 (
            .O(N__28252),
            .I(N__28241));
    LocalMux I__5833 (
            .O(N__28249),
            .I(N__28241));
    Span4Mux_h I__5832 (
            .O(N__28246),
            .I(N__28236));
    Span4Mux_h I__5831 (
            .O(N__28241),
            .I(N__28236));
    Odrv4 I__5830 (
            .O(N__28236),
            .I(dataRead3_6));
    InMux I__5829 (
            .O(N__28233),
            .I(N__28230));
    LocalMux I__5828 (
            .O(N__28230),
            .I(OutReg_0_4_i_m3_ns_1_6));
    InMux I__5827 (
            .O(N__28227),
            .I(N__28223));
    CascadeMux I__5826 (
            .O(N__28226),
            .I(N__28219));
    LocalMux I__5825 (
            .O(N__28223),
            .I(N__28216));
    CascadeMux I__5824 (
            .O(N__28222),
            .I(N__28213));
    InMux I__5823 (
            .O(N__28219),
            .I(N__28210));
    Span4Mux_h I__5822 (
            .O(N__28216),
            .I(N__28207));
    InMux I__5821 (
            .O(N__28213),
            .I(N__28204));
    LocalMux I__5820 (
            .O(N__28210),
            .I(N__28201));
    Span4Mux_h I__5819 (
            .O(N__28207),
            .I(N__28198));
    LocalMux I__5818 (
            .O(N__28204),
            .I(dataRead5_14));
    Odrv4 I__5817 (
            .O(N__28201),
            .I(dataRead5_14));
    Odrv4 I__5816 (
            .O(N__28198),
            .I(dataRead5_14));
    InMux I__5815 (
            .O(N__28191),
            .I(N__28186));
    InMux I__5814 (
            .O(N__28190),
            .I(N__28183));
    CascadeMux I__5813 (
            .O(N__28189),
            .I(N__28180));
    LocalMux I__5812 (
            .O(N__28186),
            .I(N__28177));
    LocalMux I__5811 (
            .O(N__28183),
            .I(N__28174));
    InMux I__5810 (
            .O(N__28180),
            .I(N__28171));
    Span4Mux_h I__5809 (
            .O(N__28177),
            .I(N__28168));
    Odrv4 I__5808 (
            .O(N__28174),
            .I(dataRead1_14));
    LocalMux I__5807 (
            .O(N__28171),
            .I(dataRead1_14));
    Odrv4 I__5806 (
            .O(N__28168),
            .I(dataRead1_14));
    CascadeMux I__5805 (
            .O(N__28161),
            .I(OutReg_0_5_i_m3_ns_1_14_cascade_));
    CascadeMux I__5804 (
            .O(N__28158),
            .I(OutReg_esr_RNO_2Z0Z_14_cascade_));
    InMux I__5803 (
            .O(N__28155),
            .I(N__28152));
    LocalMux I__5802 (
            .O(N__28152),
            .I(N__28149));
    Odrv12 I__5801 (
            .O(N__28149),
            .I(OutReg_esr_RNO_1Z0Z_14));
    InMux I__5800 (
            .O(N__28146),
            .I(N__28143));
    LocalMux I__5799 (
            .O(N__28143),
            .I(OutReg_esr_RNO_0Z0Z_14));
    CascadeMux I__5798 (
            .O(N__28140),
            .I(N__28134));
    CascadeMux I__5797 (
            .O(N__28139),
            .I(N__28129));
    InMux I__5796 (
            .O(N__28138),
            .I(N__28123));
    InMux I__5795 (
            .O(N__28137),
            .I(N__28118));
    InMux I__5794 (
            .O(N__28134),
            .I(N__28118));
    CascadeMux I__5793 (
            .O(N__28133),
            .I(N__28115));
    InMux I__5792 (
            .O(N__28132),
            .I(N__28112));
    InMux I__5791 (
            .O(N__28129),
            .I(N__28109));
    InMux I__5790 (
            .O(N__28128),
            .I(N__28106));
    InMux I__5789 (
            .O(N__28127),
            .I(N__28103));
    InMux I__5788 (
            .O(N__28126),
            .I(N__28098));
    LocalMux I__5787 (
            .O(N__28123),
            .I(N__28095));
    LocalMux I__5786 (
            .O(N__28118),
            .I(N__28092));
    InMux I__5785 (
            .O(N__28115),
            .I(N__28089));
    LocalMux I__5784 (
            .O(N__28112),
            .I(N__28084));
    LocalMux I__5783 (
            .O(N__28109),
            .I(N__28084));
    LocalMux I__5782 (
            .O(N__28106),
            .I(N__28081));
    LocalMux I__5781 (
            .O(N__28103),
            .I(N__28078));
    InMux I__5780 (
            .O(N__28102),
            .I(N__28075));
    InMux I__5779 (
            .O(N__28101),
            .I(N__28072));
    LocalMux I__5778 (
            .O(N__28098),
            .I(N__28067));
    Span4Mux_v I__5777 (
            .O(N__28095),
            .I(N__28067));
    Span4Mux_v I__5776 (
            .O(N__28092),
            .I(N__28062));
    LocalMux I__5775 (
            .O(N__28089),
            .I(N__28062));
    Span12Mux_s7_v I__5774 (
            .O(N__28084),
            .I(N__28059));
    Odrv4 I__5773 (
            .O(N__28081),
            .I(data_received_2_repZ0Z1));
    Odrv4 I__5772 (
            .O(N__28078),
            .I(data_received_2_repZ0Z1));
    LocalMux I__5771 (
            .O(N__28075),
            .I(data_received_2_repZ0Z1));
    LocalMux I__5770 (
            .O(N__28072),
            .I(data_received_2_repZ0Z1));
    Odrv4 I__5769 (
            .O(N__28067),
            .I(data_received_2_repZ0Z1));
    Odrv4 I__5768 (
            .O(N__28062),
            .I(data_received_2_repZ0Z1));
    Odrv12 I__5767 (
            .O(N__28059),
            .I(data_received_2_repZ0Z1));
    InMux I__5766 (
            .O(N__28044),
            .I(N__28039));
    InMux I__5765 (
            .O(N__28043),
            .I(N__28036));
    CascadeMux I__5764 (
            .O(N__28042),
            .I(N__28033));
    LocalMux I__5763 (
            .O(N__28039),
            .I(N__28028));
    LocalMux I__5762 (
            .O(N__28036),
            .I(N__28028));
    InMux I__5761 (
            .O(N__28033),
            .I(N__28025));
    Span4Mux_v I__5760 (
            .O(N__28028),
            .I(N__28022));
    LocalMux I__5759 (
            .O(N__28025),
            .I(dataRead4_3));
    Odrv4 I__5758 (
            .O(N__28022),
            .I(dataRead4_3));
    CascadeMux I__5757 (
            .O(N__28017),
            .I(N__28009));
    CascadeMux I__5756 (
            .O(N__28016),
            .I(N__28005));
    InMux I__5755 (
            .O(N__28015),
            .I(N__28000));
    InMux I__5754 (
            .O(N__28014),
            .I(N__28000));
    InMux I__5753 (
            .O(N__28013),
            .I(N__27997));
    InMux I__5752 (
            .O(N__28012),
            .I(N__27993));
    InMux I__5751 (
            .O(N__28009),
            .I(N__27990));
    InMux I__5750 (
            .O(N__28008),
            .I(N__27986));
    InMux I__5749 (
            .O(N__28005),
            .I(N__27983));
    LocalMux I__5748 (
            .O(N__28000),
            .I(N__27978));
    LocalMux I__5747 (
            .O(N__27997),
            .I(N__27978));
    CascadeMux I__5746 (
            .O(N__27996),
            .I(N__27973));
    LocalMux I__5745 (
            .O(N__27993),
            .I(N__27970));
    LocalMux I__5744 (
            .O(N__27990),
            .I(N__27967));
    InMux I__5743 (
            .O(N__27989),
            .I(N__27964));
    LocalMux I__5742 (
            .O(N__27986),
            .I(N__27961));
    LocalMux I__5741 (
            .O(N__27983),
            .I(N__27958));
    Span4Mux_v I__5740 (
            .O(N__27978),
            .I(N__27955));
    InMux I__5739 (
            .O(N__27977),
            .I(N__27952));
    InMux I__5738 (
            .O(N__27976),
            .I(N__27949));
    InMux I__5737 (
            .O(N__27973),
            .I(N__27946));
    Span4Mux_v I__5736 (
            .O(N__27970),
            .I(N__27941));
    Span4Mux_v I__5735 (
            .O(N__27967),
            .I(N__27941));
    LocalMux I__5734 (
            .O(N__27964),
            .I(N__27936));
    Span4Mux_s2_v I__5733 (
            .O(N__27961),
            .I(N__27936));
    Span4Mux_v I__5732 (
            .O(N__27958),
            .I(N__27931));
    Span4Mux_h I__5731 (
            .O(N__27955),
            .I(N__27931));
    LocalMux I__5730 (
            .O(N__27952),
            .I(data_received_0_repZ0Z1));
    LocalMux I__5729 (
            .O(N__27949),
            .I(data_received_0_repZ0Z1));
    LocalMux I__5728 (
            .O(N__27946),
            .I(data_received_0_repZ0Z1));
    Odrv4 I__5727 (
            .O(N__27941),
            .I(data_received_0_repZ0Z1));
    Odrv4 I__5726 (
            .O(N__27936),
            .I(data_received_0_repZ0Z1));
    Odrv4 I__5725 (
            .O(N__27931),
            .I(data_received_0_repZ0Z1));
    InMux I__5724 (
            .O(N__27918),
            .I(N__27914));
    InMux I__5723 (
            .O(N__27917),
            .I(N__27910));
    LocalMux I__5722 (
            .O(N__27914),
            .I(N__27907));
    InMux I__5721 (
            .O(N__27913),
            .I(N__27904));
    LocalMux I__5720 (
            .O(N__27910),
            .I(N__27901));
    Span4Mux_h I__5719 (
            .O(N__27907),
            .I(N__27898));
    LocalMux I__5718 (
            .O(N__27904),
            .I(N__27895));
    Span4Mux_v I__5717 (
            .O(N__27901),
            .I(N__27892));
    Span4Mux_v I__5716 (
            .O(N__27898),
            .I(N__27889));
    Span4Mux_h I__5715 (
            .O(N__27895),
            .I(N__27884));
    Span4Mux_h I__5714 (
            .O(N__27892),
            .I(N__27884));
    Odrv4 I__5713 (
            .O(N__27889),
            .I(dataRead5_3));
    Odrv4 I__5712 (
            .O(N__27884),
            .I(dataRead5_3));
    InMux I__5711 (
            .O(N__27879),
            .I(N__27875));
    InMux I__5710 (
            .O(N__27878),
            .I(N__27871));
    LocalMux I__5709 (
            .O(N__27875),
            .I(N__27868));
    InMux I__5708 (
            .O(N__27874),
            .I(N__27865));
    LocalMux I__5707 (
            .O(N__27871),
            .I(N__27860));
    Span4Mux_h I__5706 (
            .O(N__27868),
            .I(N__27860));
    LocalMux I__5705 (
            .O(N__27865),
            .I(N__27857));
    Span4Mux_v I__5704 (
            .O(N__27860),
            .I(N__27854));
    Span4Mux_h I__5703 (
            .O(N__27857),
            .I(N__27851));
    Odrv4 I__5702 (
            .O(N__27854),
            .I(dataRead1_3));
    Odrv4 I__5701 (
            .O(N__27851),
            .I(dataRead1_3));
    CascadeMux I__5700 (
            .O(N__27846),
            .I(OutReg_0_5_i_m3_ns_1_3_cascade_));
    InMux I__5699 (
            .O(N__27843),
            .I(N__27838));
    InMux I__5698 (
            .O(N__27842),
            .I(N__27835));
    InMux I__5697 (
            .O(N__27841),
            .I(N__27832));
    LocalMux I__5696 (
            .O(N__27838),
            .I(N__27829));
    LocalMux I__5695 (
            .O(N__27835),
            .I(N__27824));
    LocalMux I__5694 (
            .O(N__27832),
            .I(N__27824));
    Span12Mux_s10_h I__5693 (
            .O(N__27829),
            .I(N__27819));
    Span12Mux_h I__5692 (
            .O(N__27824),
            .I(N__27819));
    Odrv12 I__5691 (
            .O(N__27819),
            .I(dataRead7_3));
    CascadeMux I__5690 (
            .O(N__27816),
            .I(N__27813));
    InMux I__5689 (
            .O(N__27813),
            .I(N__27809));
    InMux I__5688 (
            .O(N__27812),
            .I(N__27806));
    LocalMux I__5687 (
            .O(N__27809),
            .I(N__27803));
    LocalMux I__5686 (
            .O(N__27806),
            .I(N__27800));
    Span4Mux_h I__5685 (
            .O(N__27803),
            .I(N__27797));
    Span4Mux_v I__5684 (
            .O(N__27800),
            .I(N__27793));
    Span4Mux_v I__5683 (
            .O(N__27797),
            .I(N__27790));
    InMux I__5682 (
            .O(N__27796),
            .I(N__27787));
    Odrv4 I__5681 (
            .O(N__27793),
            .I(dataRead6_3));
    Odrv4 I__5680 (
            .O(N__27790),
            .I(dataRead6_3));
    LocalMux I__5679 (
            .O(N__27787),
            .I(dataRead6_3));
    InMux I__5678 (
            .O(N__27780),
            .I(N__27777));
    LocalMux I__5677 (
            .O(N__27777),
            .I(N__27774));
    Odrv4 I__5676 (
            .O(N__27774),
            .I(OutReg_0_4_i_m3_ns_1_3));
    CascadeMux I__5675 (
            .O(N__27771),
            .I(OutReg_ess_RNO_1Z0Z_3_cascade_));
    InMux I__5674 (
            .O(N__27768),
            .I(N__27765));
    LocalMux I__5673 (
            .O(N__27765),
            .I(OutReg_ess_RNO_2Z0Z_3));
    CascadeMux I__5672 (
            .O(N__27762),
            .I(OutReg_ess_RNO_0Z0Z_3_cascade_));
    InMux I__5671 (
            .O(N__27759),
            .I(N__27756));
    LocalMux I__5670 (
            .O(N__27756),
            .I(OutRegZ0Z_3));
    InMux I__5669 (
            .O(N__27753),
            .I(N__27750));
    LocalMux I__5668 (
            .O(N__27750),
            .I(N__27747));
    Span4Mux_v I__5667 (
            .O(N__27747),
            .I(N__27744));
    Odrv4 I__5666 (
            .O(N__27744),
            .I(OutReg_ess_RNO_0Z0Z_4));
    InMux I__5665 (
            .O(N__27741),
            .I(N__27737));
    InMux I__5664 (
            .O(N__27740),
            .I(N__27734));
    LocalMux I__5663 (
            .O(N__27737),
            .I(N__27731));
    LocalMux I__5662 (
            .O(N__27734),
            .I(N__27728));
    Span4Mux_h I__5661 (
            .O(N__27731),
            .I(N__27725));
    Span4Mux_v I__5660 (
            .O(N__27728),
            .I(N__27721));
    Span4Mux_v I__5659 (
            .O(N__27725),
            .I(N__27718));
    InMux I__5658 (
            .O(N__27724),
            .I(N__27715));
    Odrv4 I__5657 (
            .O(N__27721),
            .I(dataRead6_6));
    Odrv4 I__5656 (
            .O(N__27718),
            .I(dataRead6_6));
    LocalMux I__5655 (
            .O(N__27715),
            .I(dataRead6_6));
    CascadeMux I__5654 (
            .O(N__27708),
            .I(N__27705));
    InMux I__5653 (
            .O(N__27705),
            .I(N__27701));
    InMux I__5652 (
            .O(N__27704),
            .I(N__27697));
    LocalMux I__5651 (
            .O(N__27701),
            .I(N__27694));
    InMux I__5650 (
            .O(N__27700),
            .I(N__27691));
    LocalMux I__5649 (
            .O(N__27697),
            .I(N__27688));
    Span4Mux_h I__5648 (
            .O(N__27694),
            .I(N__27685));
    LocalMux I__5647 (
            .O(N__27691),
            .I(N__27682));
    Span4Mux_v I__5646 (
            .O(N__27688),
            .I(N__27679));
    Span4Mux_v I__5645 (
            .O(N__27685),
            .I(N__27674));
    Span4Mux_v I__5644 (
            .O(N__27682),
            .I(N__27674));
    Odrv4 I__5643 (
            .O(N__27679),
            .I(dataRead7_6));
    Odrv4 I__5642 (
            .O(N__27674),
            .I(dataRead7_6));
    InMux I__5641 (
            .O(N__27669),
            .I(N__27666));
    LocalMux I__5640 (
            .O(N__27666),
            .I(N__27663));
    Span4Mux_v I__5639 (
            .O(N__27663),
            .I(N__27660));
    Odrv4 I__5638 (
            .O(N__27660),
            .I(OutReg_0_5_i_m3_ns_1_7));
    InMux I__5637 (
            .O(N__27657),
            .I(N__27654));
    LocalMux I__5636 (
            .O(N__27654),
            .I(N__27651));
    Odrv4 I__5635 (
            .O(N__27651),
            .I(\QuadInstance4.Quad_RNO_0_4_7 ));
    InMux I__5634 (
            .O(N__27648),
            .I(N__27645));
    LocalMux I__5633 (
            .O(N__27645),
            .I(N__27641));
    InMux I__5632 (
            .O(N__27644),
            .I(N__27637));
    Span4Mux_h I__5631 (
            .O(N__27641),
            .I(N__27634));
    InMux I__5630 (
            .O(N__27640),
            .I(N__27631));
    LocalMux I__5629 (
            .O(N__27637),
            .I(dataRead4_7));
    Odrv4 I__5628 (
            .O(N__27634),
            .I(dataRead4_7));
    LocalMux I__5627 (
            .O(N__27631),
            .I(dataRead4_7));
    InMux I__5626 (
            .O(N__27624),
            .I(N__27621));
    LocalMux I__5625 (
            .O(N__27621),
            .I(N__27618));
    Span4Mux_v I__5624 (
            .O(N__27618),
            .I(N__27615));
    Odrv4 I__5623 (
            .O(N__27615),
            .I(OutReg_0_5_i_m3_ns_1_12));
    InMux I__5622 (
            .O(N__27612),
            .I(N__27609));
    LocalMux I__5621 (
            .O(N__27609),
            .I(N__27606));
    Odrv4 I__5620 (
            .O(N__27606),
            .I(\QuadInstance4.Quad_RNO_0_4_12 ));
    CascadeMux I__5619 (
            .O(N__27603),
            .I(N__27600));
    InMux I__5618 (
            .O(N__27600),
            .I(N__27596));
    InMux I__5617 (
            .O(N__27599),
            .I(N__27592));
    LocalMux I__5616 (
            .O(N__27596),
            .I(N__27589));
    CascadeMux I__5615 (
            .O(N__27595),
            .I(N__27586));
    LocalMux I__5614 (
            .O(N__27592),
            .I(N__27583));
    Span4Mux_h I__5613 (
            .O(N__27589),
            .I(N__27580));
    InMux I__5612 (
            .O(N__27586),
            .I(N__27577));
    Odrv12 I__5611 (
            .O(N__27583),
            .I(dataRead4_12));
    Odrv4 I__5610 (
            .O(N__27580),
            .I(dataRead4_12));
    LocalMux I__5609 (
            .O(N__27577),
            .I(dataRead4_12));
    InMux I__5608 (
            .O(N__27570),
            .I(N__27566));
    InMux I__5607 (
            .O(N__27569),
            .I(N__27562));
    LocalMux I__5606 (
            .O(N__27566),
            .I(N__27559));
    InMux I__5605 (
            .O(N__27565),
            .I(N__27556));
    LocalMux I__5604 (
            .O(N__27562),
            .I(N__27553));
    Span4Mux_v I__5603 (
            .O(N__27559),
            .I(N__27548));
    LocalMux I__5602 (
            .O(N__27556),
            .I(N__27548));
    Odrv12 I__5601 (
            .O(N__27553),
            .I(dataRead4_13));
    Odrv4 I__5600 (
            .O(N__27548),
            .I(dataRead4_13));
    InMux I__5599 (
            .O(N__27543),
            .I(N__27540));
    LocalMux I__5598 (
            .O(N__27540),
            .I(N__27537));
    Span4Mux_h I__5597 (
            .O(N__27537),
            .I(N__27534));
    Span4Mux_h I__5596 (
            .O(N__27534),
            .I(N__27531));
    Odrv4 I__5595 (
            .O(N__27531),
            .I(OutReg_0_5_i_m3_ns_1_13));
    InMux I__5594 (
            .O(N__27528),
            .I(N__27524));
    InMux I__5593 (
            .O(N__27527),
            .I(N__27521));
    LocalMux I__5592 (
            .O(N__27524),
            .I(N__27518));
    LocalMux I__5591 (
            .O(N__27521),
            .I(N__27514));
    Span4Mux_v I__5590 (
            .O(N__27518),
            .I(N__27511));
    InMux I__5589 (
            .O(N__27517),
            .I(N__27508));
    Odrv4 I__5588 (
            .O(N__27514),
            .I(dataRead4_4));
    Odrv4 I__5587 (
            .O(N__27511),
            .I(dataRead4_4));
    LocalMux I__5586 (
            .O(N__27508),
            .I(dataRead4_4));
    CascadeMux I__5585 (
            .O(N__27501),
            .I(\QuadInstance4.un1_count_enable_i_a2_0_1_cascade_ ));
    CascadeMux I__5584 (
            .O(N__27498),
            .I(N__27495));
    InMux I__5583 (
            .O(N__27495),
            .I(N__27492));
    LocalMux I__5582 (
            .O(N__27492),
            .I(N__27489));
    Odrv4 I__5581 (
            .O(N__27489),
            .I(\QuadInstance4.Quad_RNIJUVR1Z0Z_4 ));
    InMux I__5580 (
            .O(N__27486),
            .I(N__27483));
    LocalMux I__5579 (
            .O(N__27483),
            .I(N__27480));
    Span4Mux_h I__5578 (
            .O(N__27480),
            .I(N__27477));
    Odrv4 I__5577 (
            .O(N__27477),
            .I(\QuadInstance4.delayedCh_AZ0Z_0 ));
    InMux I__5576 (
            .O(N__27474),
            .I(N__27469));
    InMux I__5575 (
            .O(N__27473),
            .I(N__27464));
    InMux I__5574 (
            .O(N__27472),
            .I(N__27464));
    LocalMux I__5573 (
            .O(N__27469),
            .I(\QuadInstance4.delayedCh_AZ0Z_1 ));
    LocalMux I__5572 (
            .O(N__27464),
            .I(\QuadInstance4.delayedCh_AZ0Z_1 ));
    InMux I__5571 (
            .O(N__27459),
            .I(N__27456));
    LocalMux I__5570 (
            .O(N__27456),
            .I(\QuadInstance4.delayedCh_AZ0Z_2 ));
    InMux I__5569 (
            .O(N__27453),
            .I(N__27446));
    InMux I__5568 (
            .O(N__27452),
            .I(N__27446));
    CascadeMux I__5567 (
            .O(N__27451),
            .I(N__27436));
    LocalMux I__5566 (
            .O(N__27446),
            .I(N__27433));
    CascadeMux I__5565 (
            .O(N__27445),
            .I(N__27428));
    CascadeMux I__5564 (
            .O(N__27444),
            .I(N__27424));
    CascadeMux I__5563 (
            .O(N__27443),
            .I(N__27419));
    CascadeMux I__5562 (
            .O(N__27442),
            .I(N__27416));
    CascadeMux I__5561 (
            .O(N__27441),
            .I(N__27412));
    CascadeMux I__5560 (
            .O(N__27440),
            .I(N__27409));
    InMux I__5559 (
            .O(N__27439),
            .I(N__27404));
    InMux I__5558 (
            .O(N__27436),
            .I(N__27404));
    Span12Mux_v I__5557 (
            .O(N__27433),
            .I(N__27401));
    InMux I__5556 (
            .O(N__27432),
            .I(N__27398));
    InMux I__5555 (
            .O(N__27431),
            .I(N__27393));
    InMux I__5554 (
            .O(N__27428),
            .I(N__27393));
    InMux I__5553 (
            .O(N__27427),
            .I(N__27386));
    InMux I__5552 (
            .O(N__27424),
            .I(N__27386));
    InMux I__5551 (
            .O(N__27423),
            .I(N__27386));
    InMux I__5550 (
            .O(N__27422),
            .I(N__27377));
    InMux I__5549 (
            .O(N__27419),
            .I(N__27377));
    InMux I__5548 (
            .O(N__27416),
            .I(N__27377));
    InMux I__5547 (
            .O(N__27415),
            .I(N__27377));
    InMux I__5546 (
            .O(N__27412),
            .I(N__27372));
    InMux I__5545 (
            .O(N__27409),
            .I(N__27372));
    LocalMux I__5544 (
            .O(N__27404),
            .I(N__27369));
    Odrv12 I__5543 (
            .O(N__27401),
            .I(\QuadInstance4.count_enable ));
    LocalMux I__5542 (
            .O(N__27398),
            .I(\QuadInstance4.count_enable ));
    LocalMux I__5541 (
            .O(N__27393),
            .I(\QuadInstance4.count_enable ));
    LocalMux I__5540 (
            .O(N__27386),
            .I(\QuadInstance4.count_enable ));
    LocalMux I__5539 (
            .O(N__27377),
            .I(\QuadInstance4.count_enable ));
    LocalMux I__5538 (
            .O(N__27372),
            .I(\QuadInstance4.count_enable ));
    Odrv4 I__5537 (
            .O(N__27369),
            .I(\QuadInstance4.count_enable ));
    InMux I__5536 (
            .O(N__27354),
            .I(N__27348));
    CascadeMux I__5535 (
            .O(N__27353),
            .I(N__27339));
    InMux I__5534 (
            .O(N__27352),
            .I(N__27333));
    InMux I__5533 (
            .O(N__27351),
            .I(N__27333));
    LocalMux I__5532 (
            .O(N__27348),
            .I(N__27327));
    InMux I__5531 (
            .O(N__27347),
            .I(N__27320));
    InMux I__5530 (
            .O(N__27346),
            .I(N__27320));
    InMux I__5529 (
            .O(N__27345),
            .I(N__27320));
    InMux I__5528 (
            .O(N__27344),
            .I(N__27313));
    InMux I__5527 (
            .O(N__27343),
            .I(N__27313));
    InMux I__5526 (
            .O(N__27342),
            .I(N__27313));
    InMux I__5525 (
            .O(N__27339),
            .I(N__27308));
    InMux I__5524 (
            .O(N__27338),
            .I(N__27308));
    LocalMux I__5523 (
            .O(N__27333),
            .I(N__27305));
    InMux I__5522 (
            .O(N__27332),
            .I(N__27298));
    InMux I__5521 (
            .O(N__27331),
            .I(N__27298));
    InMux I__5520 (
            .O(N__27330),
            .I(N__27298));
    Odrv12 I__5519 (
            .O(N__27327),
            .I(\QuadInstance4.un1_count_enable_i_a2_0_1 ));
    LocalMux I__5518 (
            .O(N__27320),
            .I(\QuadInstance4.un1_count_enable_i_a2_0_1 ));
    LocalMux I__5517 (
            .O(N__27313),
            .I(\QuadInstance4.un1_count_enable_i_a2_0_1 ));
    LocalMux I__5516 (
            .O(N__27308),
            .I(\QuadInstance4.un1_count_enable_i_a2_0_1 ));
    Odrv4 I__5515 (
            .O(N__27305),
            .I(\QuadInstance4.un1_count_enable_i_a2_0_1 ));
    LocalMux I__5514 (
            .O(N__27298),
            .I(\QuadInstance4.un1_count_enable_i_a2_0_1 ));
    CascadeMux I__5513 (
            .O(N__27285),
            .I(N__27282));
    InMux I__5512 (
            .O(N__27282),
            .I(N__27279));
    LocalMux I__5511 (
            .O(N__27279),
            .I(\QuadInstance4.Quad_RNIN20S1Z0Z_8 ));
    CascadeMux I__5510 (
            .O(N__27276),
            .I(N__27273));
    InMux I__5509 (
            .O(N__27273),
            .I(N__27270));
    LocalMux I__5508 (
            .O(N__27270),
            .I(N__27267));
    Odrv4 I__5507 (
            .O(N__27267),
            .I(\QuadInstance4.Quad_RNO_0_4_8 ));
    InMux I__5506 (
            .O(N__27264),
            .I(N__27260));
    InMux I__5505 (
            .O(N__27263),
            .I(N__27256));
    LocalMux I__5504 (
            .O(N__27260),
            .I(N__27253));
    CascadeMux I__5503 (
            .O(N__27259),
            .I(N__27250));
    LocalMux I__5502 (
            .O(N__27256),
            .I(N__27247));
    Span4Mux_v I__5501 (
            .O(N__27253),
            .I(N__27244));
    InMux I__5500 (
            .O(N__27250),
            .I(N__27241));
    Odrv12 I__5499 (
            .O(N__27247),
            .I(dataRead4_8));
    Odrv4 I__5498 (
            .O(N__27244),
            .I(dataRead4_8));
    LocalMux I__5497 (
            .O(N__27241),
            .I(dataRead4_8));
    CascadeMux I__5496 (
            .O(N__27234),
            .I(\QuadInstance4.count_enable_cascade_ ));
    CascadeMux I__5495 (
            .O(N__27231),
            .I(N__27228));
    InMux I__5494 (
            .O(N__27228),
            .I(N__27225));
    LocalMux I__5493 (
            .O(N__27225),
            .I(\QuadInstance4.Quad_RNIHSVR1Z0Z_2 ));
    InMux I__5492 (
            .O(N__27222),
            .I(N__27217));
    InMux I__5491 (
            .O(N__27221),
            .I(N__27214));
    InMux I__5490 (
            .O(N__27220),
            .I(N__27211));
    LocalMux I__5489 (
            .O(N__27217),
            .I(N__27206));
    LocalMux I__5488 (
            .O(N__27214),
            .I(N__27206));
    LocalMux I__5487 (
            .O(N__27211),
            .I(N__27203));
    Span4Mux_v I__5486 (
            .O(N__27206),
            .I(N__27200));
    Odrv4 I__5485 (
            .O(N__27203),
            .I(dataRead4_1));
    Odrv4 I__5484 (
            .O(N__27200),
            .I(dataRead4_1));
    CascadeMux I__5483 (
            .O(N__27195),
            .I(N__27192));
    InMux I__5482 (
            .O(N__27192),
            .I(N__27189));
    LocalMux I__5481 (
            .O(N__27189),
            .I(\QuadInstance4.Quad_RNIGRVR1Z0Z_1 ));
    InMux I__5480 (
            .O(N__27186),
            .I(N__27183));
    LocalMux I__5479 (
            .O(N__27183),
            .I(\QuadInstance4.Quad_RNO_0_4_2 ));
    CascadeMux I__5478 (
            .O(N__27180),
            .I(N__27175));
    InMux I__5477 (
            .O(N__27179),
            .I(N__27172));
    InMux I__5476 (
            .O(N__27178),
            .I(N__27169));
    InMux I__5475 (
            .O(N__27175),
            .I(N__27166));
    LocalMux I__5474 (
            .O(N__27172),
            .I(dataRead4_2));
    LocalMux I__5473 (
            .O(N__27169),
            .I(dataRead4_2));
    LocalMux I__5472 (
            .O(N__27166),
            .I(dataRead4_2));
    CascadeMux I__5471 (
            .O(N__27159),
            .I(N__27156));
    InMux I__5470 (
            .O(N__27156),
            .I(N__27153));
    LocalMux I__5469 (
            .O(N__27153),
            .I(\QuadInstance4.Quad_RNIITVR1Z0Z_3 ));
    CascadeMux I__5468 (
            .O(N__27150),
            .I(N__27147));
    InMux I__5467 (
            .O(N__27147),
            .I(N__27144));
    LocalMux I__5466 (
            .O(N__27144),
            .I(\QuadInstance4.Quad_RNI39TL1Z0Z_13 ));
    InMux I__5465 (
            .O(N__27141),
            .I(N__27138));
    LocalMux I__5464 (
            .O(N__27138),
            .I(\QuadInstance4.Quad_RNI4ATL1Z0Z_14 ));
    CascadeMux I__5463 (
            .O(N__27135),
            .I(N__27131));
    InMux I__5462 (
            .O(N__27134),
            .I(N__27128));
    InMux I__5461 (
            .O(N__27131),
            .I(N__27125));
    LocalMux I__5460 (
            .O(N__27128),
            .I(\QuadInstance4.delayedCh_BZ0Z_2 ));
    LocalMux I__5459 (
            .O(N__27125),
            .I(\QuadInstance4.delayedCh_BZ0Z_2 ));
    InMux I__5458 (
            .O(N__27120),
            .I(N__27117));
    LocalMux I__5457 (
            .O(N__27117),
            .I(N__27114));
    IoSpan4Mux I__5456 (
            .O(N__27114),
            .I(N__27111));
    Odrv4 I__5455 (
            .O(N__27111),
            .I(ch6_B_c));
    InMux I__5454 (
            .O(N__27108),
            .I(N__27105));
    LocalMux I__5453 (
            .O(N__27105),
            .I(N__27102));
    Span4Mux_h I__5452 (
            .O(N__27102),
            .I(N__27099));
    Span4Mux_v I__5451 (
            .O(N__27099),
            .I(N__27096));
    Span4Mux_v I__5450 (
            .O(N__27096),
            .I(N__27093));
    Odrv4 I__5449 (
            .O(N__27093),
            .I(\QuadInstance6.delayedCh_BZ0Z_0 ));
    IoInMux I__5448 (
            .O(N__27090),
            .I(N__27087));
    LocalMux I__5447 (
            .O(N__27087),
            .I(PWM4_obufLegalizeSB_DFFNet));
    InMux I__5446 (
            .O(N__27084),
            .I(N__27081));
    LocalMux I__5445 (
            .O(N__27081),
            .I(N__27078));
    Span4Mux_h I__5444 (
            .O(N__27078),
            .I(N__27075));
    Odrv4 I__5443 (
            .O(N__27075),
            .I(ch1_B_c));
    InMux I__5442 (
            .O(N__27072),
            .I(N__27069));
    LocalMux I__5441 (
            .O(N__27069),
            .I(N__27066));
    Span4Mux_v I__5440 (
            .O(N__27066),
            .I(N__27063));
    Odrv4 I__5439 (
            .O(N__27063),
            .I(\QuadInstance1.delayedCh_BZ0Z_0 ));
    InMux I__5438 (
            .O(N__27060),
            .I(N__27057));
    LocalMux I__5437 (
            .O(N__27057),
            .I(\QuadInstance4.Quad_RNO_0_4_5 ));
    InMux I__5436 (
            .O(N__27054),
            .I(N__27049));
    InMux I__5435 (
            .O(N__27053),
            .I(N__27046));
    InMux I__5434 (
            .O(N__27052),
            .I(N__27043));
    LocalMux I__5433 (
            .O(N__27049),
            .I(dataRead4_5));
    LocalMux I__5432 (
            .O(N__27046),
            .I(dataRead4_5));
    LocalMux I__5431 (
            .O(N__27043),
            .I(dataRead4_5));
    CascadeMux I__5430 (
            .O(N__27036),
            .I(N__27033));
    InMux I__5429 (
            .O(N__27033),
            .I(N__27030));
    LocalMux I__5428 (
            .O(N__27030),
            .I(\QuadInstance4.Quad_RNIKVVR1Z0Z_5 ));
    InMux I__5427 (
            .O(N__27027),
            .I(N__27024));
    LocalMux I__5426 (
            .O(N__27024),
            .I(\QuadInstance4.Quad_RNI28TL1Z0Z_12 ));
    InMux I__5425 (
            .O(N__27021),
            .I(N__27018));
    LocalMux I__5424 (
            .O(N__27018),
            .I(N__27015));
    Span12Mux_v I__5423 (
            .O(N__27015),
            .I(N__27012));
    Odrv12 I__5422 (
            .O(N__27012),
            .I(\PWMInstance4.un1_periodCounter12_1_0_a2_0 ));
    InMux I__5421 (
            .O(N__27009),
            .I(N__27004));
    InMux I__5420 (
            .O(N__27008),
            .I(N__26999));
    InMux I__5419 (
            .O(N__27007),
            .I(N__26999));
    LocalMux I__5418 (
            .O(N__27004),
            .I(\PWMInstance4.periodCounterZ0Z_16 ));
    LocalMux I__5417 (
            .O(N__26999),
            .I(\PWMInstance4.periodCounterZ0Z_16 ));
    InMux I__5416 (
            .O(N__26994),
            .I(N__26989));
    InMux I__5415 (
            .O(N__26993),
            .I(N__26986));
    InMux I__5414 (
            .O(N__26992),
            .I(N__26983));
    LocalMux I__5413 (
            .O(N__26989),
            .I(\PWMInstance4.periodCounterZ0Z_7 ));
    LocalMux I__5412 (
            .O(N__26986),
            .I(\PWMInstance4.periodCounterZ0Z_7 ));
    LocalMux I__5411 (
            .O(N__26983),
            .I(\PWMInstance4.periodCounterZ0Z_7 ));
    InMux I__5410 (
            .O(N__26976),
            .I(N__26967));
    InMux I__5409 (
            .O(N__26975),
            .I(N__26967));
    InMux I__5408 (
            .O(N__26974),
            .I(N__26967));
    LocalMux I__5407 (
            .O(N__26967),
            .I(N__26964));
    Span12Mux_s9_v I__5406 (
            .O(N__26964),
            .I(N__26961));
    Odrv12 I__5405 (
            .O(N__26961),
            .I(pwmWriteZ0Z_4));
    CEMux I__5404 (
            .O(N__26958),
            .I(N__26955));
    LocalMux I__5403 (
            .O(N__26955),
            .I(N__26949));
    CEMux I__5402 (
            .O(N__26954),
            .I(N__26946));
    CEMux I__5401 (
            .O(N__26953),
            .I(N__26943));
    CEMux I__5400 (
            .O(N__26952),
            .I(N__26940));
    Span4Mux_h I__5399 (
            .O(N__26949),
            .I(N__26935));
    LocalMux I__5398 (
            .O(N__26946),
            .I(N__26935));
    LocalMux I__5397 (
            .O(N__26943),
            .I(N__26931));
    LocalMux I__5396 (
            .O(N__26940),
            .I(N__26928));
    Span4Mux_v I__5395 (
            .O(N__26935),
            .I(N__26925));
    CEMux I__5394 (
            .O(N__26934),
            .I(N__26922));
    Span4Mux_h I__5393 (
            .O(N__26931),
            .I(N__26919));
    Span4Mux_h I__5392 (
            .O(N__26928),
            .I(N__26916));
    Sp12to4 I__5391 (
            .O(N__26925),
            .I(N__26911));
    LocalMux I__5390 (
            .O(N__26922),
            .I(N__26911));
    Odrv4 I__5389 (
            .O(N__26919),
            .I(\PWMInstance4.pwmWrite_0_4 ));
    Odrv4 I__5388 (
            .O(N__26916),
            .I(\PWMInstance4.pwmWrite_0_4 ));
    Odrv12 I__5387 (
            .O(N__26911),
            .I(\PWMInstance4.pwmWrite_0_4 ));
    InMux I__5386 (
            .O(N__26904),
            .I(N__26898));
    InMux I__5385 (
            .O(N__26903),
            .I(N__26898));
    LocalMux I__5384 (
            .O(N__26898),
            .I(N__26895));
    Span12Mux_s10_v I__5383 (
            .O(N__26895),
            .I(N__26892));
    Odrv12 I__5382 (
            .O(N__26892),
            .I(pwmWrite_fastZ0Z_4));
    CascadeMux I__5381 (
            .O(N__26889),
            .I(N__26884));
    InMux I__5380 (
            .O(N__26888),
            .I(N__26874));
    InMux I__5379 (
            .O(N__26887),
            .I(N__26874));
    InMux I__5378 (
            .O(N__26884),
            .I(N__26874));
    InMux I__5377 (
            .O(N__26883),
            .I(N__26874));
    LocalMux I__5376 (
            .O(N__26874),
            .I(\PWMInstance4.clkCountZ0Z_1 ));
    InMux I__5375 (
            .O(N__26871),
            .I(N__26859));
    InMux I__5374 (
            .O(N__26870),
            .I(N__26859));
    InMux I__5373 (
            .O(N__26869),
            .I(N__26859));
    InMux I__5372 (
            .O(N__26868),
            .I(N__26859));
    LocalMux I__5371 (
            .O(N__26859),
            .I(\PWMInstance4.clkCountZ0Z_0 ));
    CascadeMux I__5370 (
            .O(N__26856),
            .I(N__26852));
    InMux I__5369 (
            .O(N__26855),
            .I(N__26849));
    InMux I__5368 (
            .O(N__26852),
            .I(N__26846));
    LocalMux I__5367 (
            .O(N__26849),
            .I(\PWMInstance4.periodCounter12 ));
    LocalMux I__5366 (
            .O(N__26846),
            .I(\PWMInstance4.periodCounter12 ));
    CascadeMux I__5365 (
            .O(N__26841),
            .I(N__26838));
    InMux I__5364 (
            .O(N__26838),
            .I(N__26835));
    LocalMux I__5363 (
            .O(N__26835),
            .I(N__26830));
    InMux I__5362 (
            .O(N__26834),
            .I(N__26827));
    InMux I__5361 (
            .O(N__26833),
            .I(N__26824));
    Span4Mux_v I__5360 (
            .O(N__26830),
            .I(N__26821));
    LocalMux I__5359 (
            .O(N__26827),
            .I(\PWMInstance4.periodCounterZ0Z_15 ));
    LocalMux I__5358 (
            .O(N__26824),
            .I(\PWMInstance4.periodCounterZ0Z_15 ));
    Odrv4 I__5357 (
            .O(N__26821),
            .I(\PWMInstance4.periodCounterZ0Z_15 ));
    CascadeMux I__5356 (
            .O(N__26814),
            .I(N__26809));
    InMux I__5355 (
            .O(N__26813),
            .I(N__26806));
    InMux I__5354 (
            .O(N__26812),
            .I(N__26803));
    InMux I__5353 (
            .O(N__26809),
            .I(N__26800));
    LocalMux I__5352 (
            .O(N__26806),
            .I(\PWMInstance4.periodCounterZ0Z_1 ));
    LocalMux I__5351 (
            .O(N__26803),
            .I(\PWMInstance4.periodCounterZ0Z_1 ));
    LocalMux I__5350 (
            .O(N__26800),
            .I(\PWMInstance4.periodCounterZ0Z_1 ));
    CascadeMux I__5349 (
            .O(N__26793),
            .I(\PWMInstance4.periodCounter12_cascade_ ));
    InMux I__5348 (
            .O(N__26790),
            .I(N__26787));
    LocalMux I__5347 (
            .O(N__26787),
            .I(\PWMInstance4.un1_periodCounter12_1_0_a2_0_6 ));
    InMux I__5346 (
            .O(N__26784),
            .I(N__26781));
    LocalMux I__5345 (
            .O(N__26781),
            .I(N__26778));
    Odrv4 I__5344 (
            .O(N__26778),
            .I(\PWMInstance4.un1_periodCounter12_1_0_a2_0_10 ));
    InMux I__5343 (
            .O(N__26775),
            .I(N__26772));
    LocalMux I__5342 (
            .O(N__26772),
            .I(\PWMInstance4.un1_periodCounter12_1_0_a2_0_9 ));
    CascadeMux I__5341 (
            .O(N__26769),
            .I(\PWMInstance4.un1_periodCounter12_1_0_a2_0_14_cascade_ ));
    InMux I__5340 (
            .O(N__26766),
            .I(N__26763));
    LocalMux I__5339 (
            .O(N__26763),
            .I(N__26760));
    Odrv4 I__5338 (
            .O(N__26760),
            .I(\PWMInstance4.un1_periodCounter12_1_0_a2_0_12 ));
    CascadeMux I__5337 (
            .O(N__26757),
            .I(N__26754));
    InMux I__5336 (
            .O(N__26754),
            .I(N__26751));
    LocalMux I__5335 (
            .O(N__26751),
            .I(N__26743));
    InMux I__5334 (
            .O(N__26750),
            .I(N__26740));
    InMux I__5333 (
            .O(N__26749),
            .I(N__26737));
    InMux I__5332 (
            .O(N__26748),
            .I(N__26732));
    InMux I__5331 (
            .O(N__26747),
            .I(N__26732));
    InMux I__5330 (
            .O(N__26746),
            .I(N__26729));
    Span12Mux_s11_v I__5329 (
            .O(N__26743),
            .I(N__26726));
    LocalMux I__5328 (
            .O(N__26740),
            .I(\PWMInstance4.out_0_sqmuxa ));
    LocalMux I__5327 (
            .O(N__26737),
            .I(\PWMInstance4.out_0_sqmuxa ));
    LocalMux I__5326 (
            .O(N__26732),
            .I(\PWMInstance4.out_0_sqmuxa ));
    LocalMux I__5325 (
            .O(N__26729),
            .I(\PWMInstance4.out_0_sqmuxa ));
    Odrv12 I__5324 (
            .O(N__26726),
            .I(\PWMInstance4.out_0_sqmuxa ));
    InMux I__5323 (
            .O(N__26715),
            .I(\PWMInstance3.un1_periodCounter_2_cry_14 ));
    InMux I__5322 (
            .O(N__26712),
            .I(bfn_15_15_0_));
    CascadeMux I__5321 (
            .O(N__26709),
            .I(N__26706));
    InMux I__5320 (
            .O(N__26706),
            .I(N__26699));
    InMux I__5319 (
            .O(N__26705),
            .I(N__26699));
    InMux I__5318 (
            .O(N__26704),
            .I(N__26696));
    LocalMux I__5317 (
            .O(N__26699),
            .I(N__26693));
    LocalMux I__5316 (
            .O(N__26696),
            .I(\PWMInstance3.periodCounterZ0Z_16 ));
    Odrv4 I__5315 (
            .O(N__26693),
            .I(\PWMInstance3.periodCounterZ0Z_16 ));
    CascadeMux I__5314 (
            .O(N__26688),
            .I(N__26685));
    InMux I__5313 (
            .O(N__26685),
            .I(N__26680));
    InMux I__5312 (
            .O(N__26684),
            .I(N__26677));
    InMux I__5311 (
            .O(N__26683),
            .I(N__26674));
    LocalMux I__5310 (
            .O(N__26680),
            .I(N__26669));
    LocalMux I__5309 (
            .O(N__26677),
            .I(N__26669));
    LocalMux I__5308 (
            .O(N__26674),
            .I(\PWMInstance4.periodCounterZ0Z_13 ));
    Odrv4 I__5307 (
            .O(N__26669),
            .I(\PWMInstance4.periodCounterZ0Z_13 ));
    InMux I__5306 (
            .O(N__26664),
            .I(N__26659));
    InMux I__5305 (
            .O(N__26663),
            .I(N__26654));
    InMux I__5304 (
            .O(N__26662),
            .I(N__26654));
    LocalMux I__5303 (
            .O(N__26659),
            .I(\PWMInstance4.periodCounterZ0Z_0 ));
    LocalMux I__5302 (
            .O(N__26654),
            .I(\PWMInstance4.periodCounterZ0Z_0 ));
    InMux I__5301 (
            .O(N__26649),
            .I(N__26646));
    LocalMux I__5300 (
            .O(N__26646),
            .I(N__26643));
    Span4Mux_v I__5299 (
            .O(N__26643),
            .I(N__26640));
    Odrv4 I__5298 (
            .O(N__26640),
            .I(\PWMInstance4.PWMPulseWidthCountZ0Z_0 ));
    InMux I__5297 (
            .O(N__26637),
            .I(N__26634));
    LocalMux I__5296 (
            .O(N__26634),
            .I(N__26631));
    Span12Mux_s4_v I__5295 (
            .O(N__26631),
            .I(N__26628));
    Odrv12 I__5294 (
            .O(N__26628),
            .I(\PWMInstance4.un1_PWMPulseWidthCount_0_I_1_c_RNO_3 ));
    InMux I__5293 (
            .O(N__26625),
            .I(N__26622));
    LocalMux I__5292 (
            .O(N__26622),
            .I(\PWMInstance4.PWMPulseWidthCountZ0Z_1 ));
    InMux I__5291 (
            .O(N__26619),
            .I(N__26614));
    InMux I__5290 (
            .O(N__26618),
            .I(N__26609));
    InMux I__5289 (
            .O(N__26617),
            .I(N__26609));
    LocalMux I__5288 (
            .O(N__26614),
            .I(\PWMInstance4.periodCounterZ0Z_6 ));
    LocalMux I__5287 (
            .O(N__26609),
            .I(\PWMInstance4.periodCounterZ0Z_6 ));
    InMux I__5286 (
            .O(N__26604),
            .I(N__26601));
    LocalMux I__5285 (
            .O(N__26601),
            .I(N__26598));
    Span12Mux_s7_v I__5284 (
            .O(N__26598),
            .I(N__26595));
    Odrv12 I__5283 (
            .O(N__26595),
            .I(\PWMInstance4.un1_PWMPulseWidthCount_0_I_27_c_RNO_3 ));
    InMux I__5282 (
            .O(N__26592),
            .I(N__26589));
    LocalMux I__5281 (
            .O(N__26589),
            .I(\PWMInstance4.PWMPulseWidthCountZ0Z_6 ));
    CascadeMux I__5280 (
            .O(N__26586),
            .I(N__26583));
    InMux I__5279 (
            .O(N__26583),
            .I(N__26580));
    LocalMux I__5278 (
            .O(N__26580),
            .I(\PWMInstance4.PWMPulseWidthCountZ0Z_7 ));
    InMux I__5277 (
            .O(N__26577),
            .I(N__26574));
    LocalMux I__5276 (
            .O(N__26574),
            .I(N__26571));
    Odrv4 I__5275 (
            .O(N__26571),
            .I(\PWMInstance4.PWMPulseWidthCountZ0Z_9 ));
    CascadeMux I__5274 (
            .O(N__26568),
            .I(N__26564));
    InMux I__5273 (
            .O(N__26567),
            .I(N__26560));
    InMux I__5272 (
            .O(N__26564),
            .I(N__26555));
    InMux I__5271 (
            .O(N__26563),
            .I(N__26555));
    LocalMux I__5270 (
            .O(N__26560),
            .I(\PWMInstance4.periodCounterZ0Z_8 ));
    LocalMux I__5269 (
            .O(N__26555),
            .I(\PWMInstance4.periodCounterZ0Z_8 ));
    InMux I__5268 (
            .O(N__26550),
            .I(N__26545));
    CascadeMux I__5267 (
            .O(N__26549),
            .I(N__26542));
    InMux I__5266 (
            .O(N__26548),
            .I(N__26539));
    LocalMux I__5265 (
            .O(N__26545),
            .I(N__26536));
    InMux I__5264 (
            .O(N__26542),
            .I(N__26533));
    LocalMux I__5263 (
            .O(N__26539),
            .I(\PWMInstance4.periodCounterZ0Z_9 ));
    Odrv4 I__5262 (
            .O(N__26536),
            .I(\PWMInstance4.periodCounterZ0Z_9 ));
    LocalMux I__5261 (
            .O(N__26533),
            .I(\PWMInstance4.periodCounterZ0Z_9 ));
    InMux I__5260 (
            .O(N__26526),
            .I(N__26523));
    LocalMux I__5259 (
            .O(N__26523),
            .I(N__26520));
    Odrv4 I__5258 (
            .O(N__26520),
            .I(\PWMInstance4.PWMPulseWidthCountZ0Z_8 ));
    InMux I__5257 (
            .O(N__26517),
            .I(N__26514));
    LocalMux I__5256 (
            .O(N__26514),
            .I(N__26511));
    Span12Mux_s10_v I__5255 (
            .O(N__26511),
            .I(N__26508));
    Odrv12 I__5254 (
            .O(N__26508),
            .I(\PWMInstance4.un1_PWMPulseWidthCount_0_I_45_c_RNO_3 ));
    InMux I__5253 (
            .O(N__26505),
            .I(\PWMInstance3.un1_periodCounter_2_cry_5 ));
    InMux I__5252 (
            .O(N__26502),
            .I(\PWMInstance3.un1_periodCounter_2_cry_6 ));
    InMux I__5251 (
            .O(N__26499),
            .I(bfn_15_14_0_));
    InMux I__5250 (
            .O(N__26496),
            .I(\PWMInstance3.un1_periodCounter_2_cry_8 ));
    InMux I__5249 (
            .O(N__26493),
            .I(N__26486));
    InMux I__5248 (
            .O(N__26492),
            .I(N__26486));
    InMux I__5247 (
            .O(N__26491),
            .I(N__26483));
    LocalMux I__5246 (
            .O(N__26486),
            .I(N__26480));
    LocalMux I__5245 (
            .O(N__26483),
            .I(\PWMInstance3.periodCounterZ0Z_10 ));
    Odrv4 I__5244 (
            .O(N__26480),
            .I(\PWMInstance3.periodCounterZ0Z_10 ));
    InMux I__5243 (
            .O(N__26475),
            .I(\PWMInstance3.un1_periodCounter_2_cry_9 ));
    InMux I__5242 (
            .O(N__26472),
            .I(\PWMInstance3.un1_periodCounter_2_cry_10 ));
    InMux I__5241 (
            .O(N__26469),
            .I(\PWMInstance3.un1_periodCounter_2_cry_11 ));
    InMux I__5240 (
            .O(N__26466),
            .I(\PWMInstance3.un1_periodCounter_2_cry_12 ));
    InMux I__5239 (
            .O(N__26463),
            .I(\PWMInstance3.un1_periodCounter_2_cry_13 ));
    CascadeMux I__5238 (
            .O(N__26460),
            .I(\PWMInstance3.un1_periodCounter12_1_0_a2_0_0_cascade_ ));
    InMux I__5237 (
            .O(N__26457),
            .I(N__26454));
    LocalMux I__5236 (
            .O(N__26454),
            .I(\PWMInstance3.un1_periodCounter12_1_0_a2_0_12 ));
    InMux I__5235 (
            .O(N__26451),
            .I(N__26448));
    LocalMux I__5234 (
            .O(N__26448),
            .I(\PWMInstance3.PWMPulseWidthCountZ0Z_4 ));
    InMux I__5233 (
            .O(N__26445),
            .I(N__26442));
    LocalMux I__5232 (
            .O(N__26442),
            .I(\PWMInstance3.PWMPulseWidthCountZ0Z_11 ));
    InMux I__5231 (
            .O(N__26439),
            .I(N__26436));
    LocalMux I__5230 (
            .O(N__26436),
            .I(\PWMInstance3.PWMPulseWidthCountZ0Z_10 ));
    CascadeMux I__5229 (
            .O(N__26433),
            .I(N__26429));
    InMux I__5228 (
            .O(N__26432),
            .I(N__26425));
    InMux I__5227 (
            .O(N__26429),
            .I(N__26422));
    InMux I__5226 (
            .O(N__26428),
            .I(N__26419));
    LocalMux I__5225 (
            .O(N__26425),
            .I(\PWMInstance3.periodCounter12 ));
    LocalMux I__5224 (
            .O(N__26422),
            .I(\PWMInstance3.periodCounter12 ));
    LocalMux I__5223 (
            .O(N__26419),
            .I(\PWMInstance3.periodCounter12 ));
    InMux I__5222 (
            .O(N__26412),
            .I(\PWMInstance3.un1_periodCounter_2_cry_0 ));
    InMux I__5221 (
            .O(N__26409),
            .I(\PWMInstance3.un1_periodCounter_2_cry_1 ));
    InMux I__5220 (
            .O(N__26406),
            .I(\PWMInstance3.un1_periodCounter_2_cry_2 ));
    InMux I__5219 (
            .O(N__26403),
            .I(N__26398));
    InMux I__5218 (
            .O(N__26402),
            .I(N__26393));
    InMux I__5217 (
            .O(N__26401),
            .I(N__26393));
    LocalMux I__5216 (
            .O(N__26398),
            .I(\PWMInstance3.periodCounterZ0Z_4 ));
    LocalMux I__5215 (
            .O(N__26393),
            .I(\PWMInstance3.periodCounterZ0Z_4 ));
    InMux I__5214 (
            .O(N__26388),
            .I(\PWMInstance3.un1_periodCounter_2_cry_3 ));
    InMux I__5213 (
            .O(N__26385),
            .I(\PWMInstance3.un1_periodCounter_2_cry_4 ));
    CascadeMux I__5212 (
            .O(N__26382),
            .I(OutReg_ess_RNO_2Z0Z_7_cascade_));
    CascadeMux I__5211 (
            .O(N__26379),
            .I(OutReg_ess_RNO_0Z0Z_7_cascade_));
    InMux I__5210 (
            .O(N__26376),
            .I(N__26371));
    InMux I__5209 (
            .O(N__26375),
            .I(N__26368));
    InMux I__5208 (
            .O(N__26374),
            .I(N__26365));
    LocalMux I__5207 (
            .O(N__26371),
            .I(N__26362));
    LocalMux I__5206 (
            .O(N__26368),
            .I(N__26359));
    LocalMux I__5205 (
            .O(N__26365),
            .I(N__26356));
    Span4Mux_h I__5204 (
            .O(N__26362),
            .I(N__26353));
    Span4Mux_h I__5203 (
            .O(N__26359),
            .I(N__26350));
    Span4Mux_h I__5202 (
            .O(N__26356),
            .I(N__26345));
    Span4Mux_v I__5201 (
            .O(N__26353),
            .I(N__26345));
    Odrv4 I__5200 (
            .O(N__26350),
            .I(dataRead2_7));
    Odrv4 I__5199 (
            .O(N__26345),
            .I(dataRead2_7));
    CascadeMux I__5198 (
            .O(N__26340),
            .I(N__26337));
    InMux I__5197 (
            .O(N__26337),
            .I(N__26333));
    InMux I__5196 (
            .O(N__26336),
            .I(N__26330));
    LocalMux I__5195 (
            .O(N__26333),
            .I(N__26326));
    LocalMux I__5194 (
            .O(N__26330),
            .I(N__26323));
    InMux I__5193 (
            .O(N__26329),
            .I(N__26320));
    Span4Mux_h I__5192 (
            .O(N__26326),
            .I(N__26317));
    Span4Mux_v I__5191 (
            .O(N__26323),
            .I(N__26312));
    LocalMux I__5190 (
            .O(N__26320),
            .I(N__26312));
    Span4Mux_v I__5189 (
            .O(N__26317),
            .I(N__26309));
    Odrv4 I__5188 (
            .O(N__26312),
            .I(dataRead3_7));
    Odrv4 I__5187 (
            .O(N__26309),
            .I(dataRead3_7));
    InMux I__5186 (
            .O(N__26304),
            .I(N__26300));
    InMux I__5185 (
            .O(N__26303),
            .I(N__26297));
    LocalMux I__5184 (
            .O(N__26300),
            .I(N__26294));
    LocalMux I__5183 (
            .O(N__26297),
            .I(N__26291));
    Span4Mux_v I__5182 (
            .O(N__26294),
            .I(N__26288));
    Span12Mux_v I__5181 (
            .O(N__26291),
            .I(N__26284));
    Span4Mux_v I__5180 (
            .O(N__26288),
            .I(N__26281));
    InMux I__5179 (
            .O(N__26287),
            .I(N__26278));
    Odrv12 I__5178 (
            .O(N__26284),
            .I(dataRead6_7));
    Odrv4 I__5177 (
            .O(N__26281),
            .I(dataRead6_7));
    LocalMux I__5176 (
            .O(N__26278),
            .I(dataRead6_7));
    InMux I__5175 (
            .O(N__26271),
            .I(N__26267));
    InMux I__5174 (
            .O(N__26270),
            .I(N__26264));
    LocalMux I__5173 (
            .O(N__26267),
            .I(N__26261));
    LocalMux I__5172 (
            .O(N__26264),
            .I(N__26258));
    Span4Mux_v I__5171 (
            .O(N__26261),
            .I(N__26252));
    Span4Mux_h I__5170 (
            .O(N__26258),
            .I(N__26252));
    InMux I__5169 (
            .O(N__26257),
            .I(N__26249));
    Span4Mux_h I__5168 (
            .O(N__26252),
            .I(N__26244));
    LocalMux I__5167 (
            .O(N__26249),
            .I(N__26244));
    Span4Mux_v I__5166 (
            .O(N__26244),
            .I(N__26241));
    Odrv4 I__5165 (
            .O(N__26241),
            .I(dataRead7_7));
    CascadeMux I__5164 (
            .O(N__26238),
            .I(OutReg_0_4_i_m3_ns_1_7_cascade_));
    InMux I__5163 (
            .O(N__26235),
            .I(N__26232));
    LocalMux I__5162 (
            .O(N__26232),
            .I(OutReg_ess_RNO_1Z0Z_7));
    InMux I__5161 (
            .O(N__26229),
            .I(N__26226));
    LocalMux I__5160 (
            .O(N__26226),
            .I(N__26223));
    Odrv4 I__5159 (
            .O(N__26223),
            .I(OutReg_ess_RNO_0Z0Z_9));
    CascadeMux I__5158 (
            .O(N__26220),
            .I(N__26217));
    InMux I__5157 (
            .O(N__26217),
            .I(N__26214));
    LocalMux I__5156 (
            .O(N__26214),
            .I(N__26211));
    Span4Mux_v I__5155 (
            .O(N__26211),
            .I(N__26208));
    Odrv4 I__5154 (
            .O(N__26208),
            .I(OutRegZ0Z_13));
    CascadeMux I__5153 (
            .O(N__26205),
            .I(N__26202));
    InMux I__5152 (
            .O(N__26202),
            .I(N__26199));
    LocalMux I__5151 (
            .O(N__26199),
            .I(N__26196));
    Span4Mux_h I__5150 (
            .O(N__26196),
            .I(N__26193));
    Odrv4 I__5149 (
            .O(N__26193),
            .I(OutRegZ0Z_14));
    InMux I__5148 (
            .O(N__26190),
            .I(N__26187));
    LocalMux I__5147 (
            .O(N__26187),
            .I(\PWMInstance3.PWMPulseWidthCountZ0Z_5 ));
    CEMux I__5146 (
            .O(N__26184),
            .I(N__26163));
    CEMux I__5145 (
            .O(N__26183),
            .I(N__26163));
    CEMux I__5144 (
            .O(N__26182),
            .I(N__26163));
    CEMux I__5143 (
            .O(N__26181),
            .I(N__26163));
    CEMux I__5142 (
            .O(N__26180),
            .I(N__26163));
    CEMux I__5141 (
            .O(N__26179),
            .I(N__26163));
    CEMux I__5140 (
            .O(N__26178),
            .I(N__26163));
    GlobalMux I__5139 (
            .O(N__26163),
            .I(N__26160));
    gio2CtrlBuf I__5138 (
            .O(N__26160),
            .I(N_45_0_g));
    SRMux I__5137 (
            .O(N__26157),
            .I(N__26136));
    SRMux I__5136 (
            .O(N__26156),
            .I(N__26136));
    SRMux I__5135 (
            .O(N__26155),
            .I(N__26136));
    SRMux I__5134 (
            .O(N__26154),
            .I(N__26136));
    SRMux I__5133 (
            .O(N__26153),
            .I(N__26136));
    SRMux I__5132 (
            .O(N__26152),
            .I(N__26136));
    SRMux I__5131 (
            .O(N__26151),
            .I(N__26136));
    GlobalMux I__5130 (
            .O(N__26136),
            .I(N__26133));
    gio2CtrlBuf I__5129 (
            .O(N__26133),
            .I(N_1187_g));
    InMux I__5128 (
            .O(N__26130),
            .I(N__26127));
    LocalMux I__5127 (
            .O(N__26127),
            .I(N__26124));
    Odrv12 I__5126 (
            .O(N__26124),
            .I(\QuadInstance4.Quad_RNO_0_4_13 ));
    InMux I__5125 (
            .O(N__26121),
            .I(N__26118));
    LocalMux I__5124 (
            .O(N__26118),
            .I(N__26115));
    Odrv12 I__5123 (
            .O(N__26115),
            .I(\QuadInstance7.Quad_RNO_0_7_13 ));
    InMux I__5122 (
            .O(N__26112),
            .I(N__26109));
    LocalMux I__5121 (
            .O(N__26109),
            .I(N__26104));
    InMux I__5120 (
            .O(N__26108),
            .I(N__26101));
    CascadeMux I__5119 (
            .O(N__26107),
            .I(N__26098));
    Span4Mux_h I__5118 (
            .O(N__26104),
            .I(N__26093));
    LocalMux I__5117 (
            .O(N__26101),
            .I(N__26093));
    InMux I__5116 (
            .O(N__26098),
            .I(N__26090));
    Span4Mux_h I__5115 (
            .O(N__26093),
            .I(N__26087));
    LocalMux I__5114 (
            .O(N__26090),
            .I(N__26084));
    Odrv4 I__5113 (
            .O(N__26087),
            .I(dataRead7_13));
    Odrv12 I__5112 (
            .O(N__26084),
            .I(dataRead7_13));
    InMux I__5111 (
            .O(N__26079),
            .I(N__26076));
    LocalMux I__5110 (
            .O(N__26076),
            .I(N__26073));
    Odrv12 I__5109 (
            .O(N__26073),
            .I(\QuadInstance4.Quad_RNO_0_4_3 ));
    InMux I__5108 (
            .O(N__26070),
            .I(N__26067));
    LocalMux I__5107 (
            .O(N__26067),
            .I(N__26064));
    Span4Mux_h I__5106 (
            .O(N__26064),
            .I(N__26061));
    Span4Mux_h I__5105 (
            .O(N__26061),
            .I(N__26058));
    Odrv4 I__5104 (
            .O(N__26058),
            .I(\QuadInstance7.Quad_RNO_0_7_3 ));
    InMux I__5103 (
            .O(N__26055),
            .I(N__26047));
    InMux I__5102 (
            .O(N__26054),
            .I(N__26047));
    InMux I__5101 (
            .O(N__26053),
            .I(N__26044));
    InMux I__5100 (
            .O(N__26052),
            .I(N__26034));
    LocalMux I__5099 (
            .O(N__26047),
            .I(N__26031));
    LocalMux I__5098 (
            .O(N__26044),
            .I(N__26028));
    InMux I__5097 (
            .O(N__26043),
            .I(N__26025));
    CascadeMux I__5096 (
            .O(N__26042),
            .I(N__26022));
    InMux I__5095 (
            .O(N__26041),
            .I(N__26015));
    InMux I__5094 (
            .O(N__26040),
            .I(N__26015));
    InMux I__5093 (
            .O(N__26039),
            .I(N__26015));
    InMux I__5092 (
            .O(N__26038),
            .I(N__26008));
    CascadeMux I__5091 (
            .O(N__26037),
            .I(N__26005));
    LocalMux I__5090 (
            .O(N__26034),
            .I(N__26001));
    Span4Mux_v I__5089 (
            .O(N__26031),
            .I(N__25994));
    Span4Mux_v I__5088 (
            .O(N__26028),
            .I(N__25994));
    LocalMux I__5087 (
            .O(N__26025),
            .I(N__25994));
    InMux I__5086 (
            .O(N__26022),
            .I(N__25991));
    LocalMux I__5085 (
            .O(N__26015),
            .I(N__25988));
    InMux I__5084 (
            .O(N__26014),
            .I(N__25983));
    InMux I__5083 (
            .O(N__26013),
            .I(N__25983));
    InMux I__5082 (
            .O(N__26012),
            .I(N__25980));
    CascadeMux I__5081 (
            .O(N__26011),
            .I(N__25977));
    LocalMux I__5080 (
            .O(N__26008),
            .I(N__25966));
    InMux I__5079 (
            .O(N__26005),
            .I(N__25961));
    InMux I__5078 (
            .O(N__26004),
            .I(N__25961));
    Span4Mux_v I__5077 (
            .O(N__26001),
            .I(N__25956));
    Span4Mux_h I__5076 (
            .O(N__25994),
            .I(N__25956));
    LocalMux I__5075 (
            .O(N__25991),
            .I(N__25951));
    Span4Mux_v I__5074 (
            .O(N__25988),
            .I(N__25951));
    LocalMux I__5073 (
            .O(N__25983),
            .I(N__25946));
    LocalMux I__5072 (
            .O(N__25980),
            .I(N__25946));
    InMux I__5071 (
            .O(N__25977),
            .I(N__25943));
    InMux I__5070 (
            .O(N__25976),
            .I(N__25936));
    InMux I__5069 (
            .O(N__25975),
            .I(N__25936));
    InMux I__5068 (
            .O(N__25974),
            .I(N__25936));
    CascadeMux I__5067 (
            .O(N__25973),
            .I(N__25932));
    CascadeMux I__5066 (
            .O(N__25972),
            .I(N__25929));
    CascadeMux I__5065 (
            .O(N__25971),
            .I(N__25924));
    CascadeMux I__5064 (
            .O(N__25970),
            .I(N__25921));
    InMux I__5063 (
            .O(N__25969),
            .I(N__25914));
    Span4Mux_h I__5062 (
            .O(N__25966),
            .I(N__25907));
    LocalMux I__5061 (
            .O(N__25961),
            .I(N__25907));
    Span4Mux_h I__5060 (
            .O(N__25956),
            .I(N__25907));
    Span4Mux_h I__5059 (
            .O(N__25951),
            .I(N__25902));
    Span4Mux_v I__5058 (
            .O(N__25946),
            .I(N__25902));
    LocalMux I__5057 (
            .O(N__25943),
            .I(N__25897));
    LocalMux I__5056 (
            .O(N__25936),
            .I(N__25897));
    InMux I__5055 (
            .O(N__25935),
            .I(N__25888));
    InMux I__5054 (
            .O(N__25932),
            .I(N__25888));
    InMux I__5053 (
            .O(N__25929),
            .I(N__25888));
    InMux I__5052 (
            .O(N__25928),
            .I(N__25888));
    InMux I__5051 (
            .O(N__25927),
            .I(N__25877));
    InMux I__5050 (
            .O(N__25924),
            .I(N__25877));
    InMux I__5049 (
            .O(N__25921),
            .I(N__25877));
    InMux I__5048 (
            .O(N__25920),
            .I(N__25877));
    InMux I__5047 (
            .O(N__25919),
            .I(N__25877));
    InMux I__5046 (
            .O(N__25918),
            .I(N__25872));
    InMux I__5045 (
            .O(N__25917),
            .I(N__25872));
    LocalMux I__5044 (
            .O(N__25914),
            .I(quadWriteZ0Z_7));
    Odrv4 I__5043 (
            .O(N__25907),
            .I(quadWriteZ0Z_7));
    Odrv4 I__5042 (
            .O(N__25902),
            .I(quadWriteZ0Z_7));
    Odrv4 I__5041 (
            .O(N__25897),
            .I(quadWriteZ0Z_7));
    LocalMux I__5040 (
            .O(N__25888),
            .I(quadWriteZ0Z_7));
    LocalMux I__5039 (
            .O(N__25877),
            .I(quadWriteZ0Z_7));
    LocalMux I__5038 (
            .O(N__25872),
            .I(quadWriteZ0Z_7));
    InMux I__5037 (
            .O(N__25857),
            .I(N__25854));
    LocalMux I__5036 (
            .O(N__25854),
            .I(N__25851));
    Span4Mux_h I__5035 (
            .O(N__25851),
            .I(N__25848));
    Span4Mux_h I__5034 (
            .O(N__25848),
            .I(N__25845));
    Odrv4 I__5033 (
            .O(N__25845),
            .I(\QuadInstance7.Quad_RNO_0_6_1 ));
    InMux I__5032 (
            .O(N__25842),
            .I(N__25838));
    InMux I__5031 (
            .O(N__25841),
            .I(N__25835));
    LocalMux I__5030 (
            .O(N__25838),
            .I(N__25831));
    LocalMux I__5029 (
            .O(N__25835),
            .I(N__25828));
    InMux I__5028 (
            .O(N__25834),
            .I(N__25825));
    Span4Mux_h I__5027 (
            .O(N__25831),
            .I(N__25822));
    Sp12to4 I__5026 (
            .O(N__25828),
            .I(N__25819));
    LocalMux I__5025 (
            .O(N__25825),
            .I(N__25816));
    Span4Mux_h I__5024 (
            .O(N__25822),
            .I(N__25813));
    Odrv12 I__5023 (
            .O(N__25819),
            .I(dataRead7_1));
    Odrv4 I__5022 (
            .O(N__25816),
            .I(dataRead7_1));
    Odrv4 I__5021 (
            .O(N__25813),
            .I(dataRead7_1));
    InMux I__5020 (
            .O(N__25806),
            .I(N__25803));
    LocalMux I__5019 (
            .O(N__25803),
            .I(N__25792));
    InMux I__5018 (
            .O(N__25802),
            .I(N__25789));
    InMux I__5017 (
            .O(N__25801),
            .I(N__25786));
    InMux I__5016 (
            .O(N__25800),
            .I(N__25779));
    InMux I__5015 (
            .O(N__25799),
            .I(N__25779));
    InMux I__5014 (
            .O(N__25798),
            .I(N__25779));
    InMux I__5013 (
            .O(N__25797),
            .I(N__25773));
    InMux I__5012 (
            .O(N__25796),
            .I(N__25773));
    InMux I__5011 (
            .O(N__25795),
            .I(N__25769));
    Span4Mux_h I__5010 (
            .O(N__25792),
            .I(N__25764));
    LocalMux I__5009 (
            .O(N__25789),
            .I(N__25764));
    LocalMux I__5008 (
            .O(N__25786),
            .I(N__25761));
    LocalMux I__5007 (
            .O(N__25779),
            .I(N__25758));
    InMux I__5006 (
            .O(N__25778),
            .I(N__25753));
    LocalMux I__5005 (
            .O(N__25773),
            .I(N__25750));
    InMux I__5004 (
            .O(N__25772),
            .I(N__25747));
    LocalMux I__5003 (
            .O(N__25769),
            .I(N__25744));
    Span4Mux_v I__5002 (
            .O(N__25764),
            .I(N__25739));
    Span4Mux_h I__5001 (
            .O(N__25761),
            .I(N__25739));
    Span4Mux_h I__5000 (
            .O(N__25758),
            .I(N__25736));
    CascadeMux I__4999 (
            .O(N__25757),
            .I(N__25717));
    InMux I__4998 (
            .O(N__25756),
            .I(N__25712));
    LocalMux I__4997 (
            .O(N__25753),
            .I(N__25707));
    Span4Mux_h I__4996 (
            .O(N__25750),
            .I(N__25707));
    LocalMux I__4995 (
            .O(N__25747),
            .I(N__25702));
    Span4Mux_v I__4994 (
            .O(N__25744),
            .I(N__25702));
    Span4Mux_h I__4993 (
            .O(N__25739),
            .I(N__25697));
    Span4Mux_h I__4992 (
            .O(N__25736),
            .I(N__25697));
    InMux I__4991 (
            .O(N__25735),
            .I(N__25680));
    InMux I__4990 (
            .O(N__25734),
            .I(N__25680));
    InMux I__4989 (
            .O(N__25733),
            .I(N__25680));
    InMux I__4988 (
            .O(N__25732),
            .I(N__25680));
    InMux I__4987 (
            .O(N__25731),
            .I(N__25680));
    InMux I__4986 (
            .O(N__25730),
            .I(N__25680));
    InMux I__4985 (
            .O(N__25729),
            .I(N__25680));
    InMux I__4984 (
            .O(N__25728),
            .I(N__25680));
    InMux I__4983 (
            .O(N__25727),
            .I(N__25669));
    InMux I__4982 (
            .O(N__25726),
            .I(N__25669));
    InMux I__4981 (
            .O(N__25725),
            .I(N__25669));
    InMux I__4980 (
            .O(N__25724),
            .I(N__25669));
    InMux I__4979 (
            .O(N__25723),
            .I(N__25669));
    InMux I__4978 (
            .O(N__25722),
            .I(N__25656));
    InMux I__4977 (
            .O(N__25721),
            .I(N__25656));
    InMux I__4976 (
            .O(N__25720),
            .I(N__25656));
    InMux I__4975 (
            .O(N__25717),
            .I(N__25656));
    InMux I__4974 (
            .O(N__25716),
            .I(N__25656));
    InMux I__4973 (
            .O(N__25715),
            .I(N__25656));
    LocalMux I__4972 (
            .O(N__25712),
            .I(quadWriteZ0Z_5));
    Odrv4 I__4971 (
            .O(N__25707),
            .I(quadWriteZ0Z_5));
    Odrv4 I__4970 (
            .O(N__25702),
            .I(quadWriteZ0Z_5));
    Odrv4 I__4969 (
            .O(N__25697),
            .I(quadWriteZ0Z_5));
    LocalMux I__4968 (
            .O(N__25680),
            .I(quadWriteZ0Z_5));
    LocalMux I__4967 (
            .O(N__25669),
            .I(quadWriteZ0Z_5));
    LocalMux I__4966 (
            .O(N__25656),
            .I(quadWriteZ0Z_5));
    InMux I__4965 (
            .O(N__25641),
            .I(N__25638));
    LocalMux I__4964 (
            .O(N__25638),
            .I(N__25635));
    Span4Mux_h I__4963 (
            .O(N__25635),
            .I(N__25632));
    Span4Mux_h I__4962 (
            .O(N__25632),
            .I(N__25629));
    Odrv4 I__4961 (
            .O(N__25629),
            .I(\QuadInstance5.Quad_RNO_0_5_3 ));
    IoInMux I__4960 (
            .O(N__25626),
            .I(N__25623));
    LocalMux I__4959 (
            .O(N__25623),
            .I(N__25620));
    Span4Mux_s3_v I__4958 (
            .O(N__25620),
            .I(N__25617));
    Span4Mux_v I__4957 (
            .O(N__25617),
            .I(N__25614));
    Span4Mux_v I__4956 (
            .O(N__25614),
            .I(N__25611));
    Odrv4 I__4955 (
            .O(N__25611),
            .I(GB_BUFFER_RST_c_i_g_THRU_CO));
    InMux I__4954 (
            .O(N__25608),
            .I(N__25604));
    InMux I__4953 (
            .O(N__25607),
            .I(N__25601));
    LocalMux I__4952 (
            .O(N__25604),
            .I(N__25598));
    LocalMux I__4951 (
            .O(N__25601),
            .I(N__25594));
    Span4Mux_h I__4950 (
            .O(N__25598),
            .I(N__25591));
    CascadeMux I__4949 (
            .O(N__25597),
            .I(N__25588));
    Span4Mux_h I__4948 (
            .O(N__25594),
            .I(N__25583));
    Span4Mux_v I__4947 (
            .O(N__25591),
            .I(N__25583));
    InMux I__4946 (
            .O(N__25588),
            .I(N__25580));
    Odrv4 I__4945 (
            .O(N__25583),
            .I(dataRead5_7));
    LocalMux I__4944 (
            .O(N__25580),
            .I(dataRead5_7));
    CascadeMux I__4943 (
            .O(N__25575),
            .I(N__25572));
    InMux I__4942 (
            .O(N__25572),
            .I(N__25569));
    LocalMux I__4941 (
            .O(N__25569),
            .I(N__25564));
    InMux I__4940 (
            .O(N__25568),
            .I(N__25561));
    InMux I__4939 (
            .O(N__25567),
            .I(N__25558));
    Span4Mux_v I__4938 (
            .O(N__25564),
            .I(N__25555));
    LocalMux I__4937 (
            .O(N__25561),
            .I(N__25550));
    LocalMux I__4936 (
            .O(N__25558),
            .I(N__25550));
    Odrv4 I__4935 (
            .O(N__25555),
            .I(dataRead1_7));
    Odrv12 I__4934 (
            .O(N__25550),
            .I(dataRead1_7));
    InMux I__4933 (
            .O(N__25545),
            .I(N__25541));
    InMux I__4932 (
            .O(N__25544),
            .I(N__25538));
    LocalMux I__4931 (
            .O(N__25541),
            .I(N__25535));
    LocalMux I__4930 (
            .O(N__25538),
            .I(N__25532));
    Span4Mux_v I__4929 (
            .O(N__25535),
            .I(N__25526));
    Span4Mux_h I__4928 (
            .O(N__25532),
            .I(N__25526));
    InMux I__4927 (
            .O(N__25531),
            .I(N__25523));
    Odrv4 I__4926 (
            .O(N__25526),
            .I(dataRead1_9));
    LocalMux I__4925 (
            .O(N__25523),
            .I(dataRead1_9));
    CascadeMux I__4924 (
            .O(N__25518),
            .I(N__25515));
    InMux I__4923 (
            .O(N__25515),
            .I(N__25511));
    InMux I__4922 (
            .O(N__25514),
            .I(N__25508));
    LocalMux I__4921 (
            .O(N__25511),
            .I(N__25504));
    LocalMux I__4920 (
            .O(N__25508),
            .I(N__25501));
    InMux I__4919 (
            .O(N__25507),
            .I(N__25498));
    Span4Mux_h I__4918 (
            .O(N__25504),
            .I(N__25495));
    Span4Mux_v I__4917 (
            .O(N__25501),
            .I(N__25490));
    LocalMux I__4916 (
            .O(N__25498),
            .I(N__25490));
    Odrv4 I__4915 (
            .O(N__25495),
            .I(dataRead5_9));
    Odrv4 I__4914 (
            .O(N__25490),
            .I(dataRead5_9));
    CascadeMux I__4913 (
            .O(N__25485),
            .I(OutReg_ess_RNO_2Z0Z_9_cascade_));
    InMux I__4912 (
            .O(N__25482),
            .I(N__25477));
    InMux I__4911 (
            .O(N__25481),
            .I(N__25474));
    InMux I__4910 (
            .O(N__25480),
            .I(N__25471));
    LocalMux I__4909 (
            .O(N__25477),
            .I(N__25468));
    LocalMux I__4908 (
            .O(N__25474),
            .I(N__25463));
    LocalMux I__4907 (
            .O(N__25471),
            .I(N__25463));
    Span4Mux_h I__4906 (
            .O(N__25468),
            .I(N__25460));
    Span4Mux_v I__4905 (
            .O(N__25463),
            .I(N__25455));
    Span4Mux_h I__4904 (
            .O(N__25460),
            .I(N__25455));
    Odrv4 I__4903 (
            .O(N__25455),
            .I(dataRead3_9));
    CascadeMux I__4902 (
            .O(N__25452),
            .I(N__25449));
    InMux I__4901 (
            .O(N__25449),
            .I(N__25446));
    LocalMux I__4900 (
            .O(N__25446),
            .I(N__25443));
    Span4Mux_v I__4899 (
            .O(N__25443),
            .I(N__25439));
    InMux I__4898 (
            .O(N__25442),
            .I(N__25435));
    Span4Mux_h I__4897 (
            .O(N__25439),
            .I(N__25432));
    InMux I__4896 (
            .O(N__25438),
            .I(N__25429));
    LocalMux I__4895 (
            .O(N__25435),
            .I(N__25424));
    Span4Mux_h I__4894 (
            .O(N__25432),
            .I(N__25424));
    LocalMux I__4893 (
            .O(N__25429),
            .I(dataRead2_9));
    Odrv4 I__4892 (
            .O(N__25424),
            .I(dataRead2_9));
    InMux I__4891 (
            .O(N__25419),
            .I(N__25415));
    InMux I__4890 (
            .O(N__25418),
            .I(N__25411));
    LocalMux I__4889 (
            .O(N__25415),
            .I(N__25408));
    InMux I__4888 (
            .O(N__25414),
            .I(N__25405));
    LocalMux I__4887 (
            .O(N__25411),
            .I(N__25400));
    Span4Mux_h I__4886 (
            .O(N__25408),
            .I(N__25400));
    LocalMux I__4885 (
            .O(N__25405),
            .I(N__25397));
    Odrv4 I__4884 (
            .O(N__25400),
            .I(dataRead6_9));
    Odrv4 I__4883 (
            .O(N__25397),
            .I(dataRead6_9));
    InMux I__4882 (
            .O(N__25392),
            .I(N__25388));
    InMux I__4881 (
            .O(N__25391),
            .I(N__25384));
    LocalMux I__4880 (
            .O(N__25388),
            .I(N__25381));
    InMux I__4879 (
            .O(N__25387),
            .I(N__25378));
    LocalMux I__4878 (
            .O(N__25384),
            .I(N__25375));
    Span4Mux_h I__4877 (
            .O(N__25381),
            .I(N__25370));
    LocalMux I__4876 (
            .O(N__25378),
            .I(N__25370));
    Span12Mux_v I__4875 (
            .O(N__25375),
            .I(N__25367));
    Span4Mux_v I__4874 (
            .O(N__25370),
            .I(N__25364));
    Odrv12 I__4873 (
            .O(N__25367),
            .I(dataRead7_9));
    Odrv4 I__4872 (
            .O(N__25364),
            .I(dataRead7_9));
    CascadeMux I__4871 (
            .O(N__25359),
            .I(OutReg_0_4_i_m3_ns_1_9_cascade_));
    InMux I__4870 (
            .O(N__25356),
            .I(N__25353));
    LocalMux I__4869 (
            .O(N__25353),
            .I(OutReg_ess_RNO_1Z0Z_9));
    CascadeMux I__4868 (
            .O(N__25350),
            .I(N__25345));
    InMux I__4867 (
            .O(N__25349),
            .I(N__25342));
    InMux I__4866 (
            .O(N__25348),
            .I(N__25339));
    InMux I__4865 (
            .O(N__25345),
            .I(N__25336));
    LocalMux I__4864 (
            .O(N__25342),
            .I(N__25331));
    LocalMux I__4863 (
            .O(N__25339),
            .I(N__25331));
    LocalMux I__4862 (
            .O(N__25336),
            .I(N__25328));
    Span4Mux_v I__4861 (
            .O(N__25331),
            .I(N__25323));
    Span4Mux_v I__4860 (
            .O(N__25328),
            .I(N__25323));
    Span4Mux_h I__4859 (
            .O(N__25323),
            .I(N__25320));
    Odrv4 I__4858 (
            .O(N__25320),
            .I(dataRead4_9));
    InMux I__4857 (
            .O(N__25317),
            .I(N__25314));
    LocalMux I__4856 (
            .O(N__25314),
            .I(OutReg_0_5_i_m3_ns_1_9));
    InMux I__4855 (
            .O(N__25311),
            .I(N__25307));
    InMux I__4854 (
            .O(N__25310),
            .I(N__25304));
    LocalMux I__4853 (
            .O(N__25307),
            .I(N__25300));
    LocalMux I__4852 (
            .O(N__25304),
            .I(N__25297));
    InMux I__4851 (
            .O(N__25303),
            .I(N__25294));
    Span4Mux_v I__4850 (
            .O(N__25300),
            .I(N__25291));
    Span4Mux_h I__4849 (
            .O(N__25297),
            .I(N__25286));
    LocalMux I__4848 (
            .O(N__25294),
            .I(N__25286));
    Odrv4 I__4847 (
            .O(N__25291),
            .I(dataRead1_6));
    Odrv4 I__4846 (
            .O(N__25286),
            .I(dataRead1_6));
    InMux I__4845 (
            .O(N__25281),
            .I(N__25277));
    InMux I__4844 (
            .O(N__25280),
            .I(N__25274));
    LocalMux I__4843 (
            .O(N__25277),
            .I(N__25271));
    LocalMux I__4842 (
            .O(N__25274),
            .I(N__25268));
    Span4Mux_h I__4841 (
            .O(N__25271),
            .I(N__25262));
    Span4Mux_h I__4840 (
            .O(N__25268),
            .I(N__25262));
    InMux I__4839 (
            .O(N__25267),
            .I(N__25259));
    Odrv4 I__4838 (
            .O(N__25262),
            .I(dataRead5_6));
    LocalMux I__4837 (
            .O(N__25259),
            .I(dataRead5_6));
    CascadeMux I__4836 (
            .O(N__25254),
            .I(OutReg_0_5_i_m3_ns_1_6_cascade_));
    CascadeMux I__4835 (
            .O(N__25251),
            .I(N__25248));
    InMux I__4834 (
            .O(N__25248),
            .I(N__25245));
    LocalMux I__4833 (
            .O(N__25245),
            .I(N__25242));
    Odrv4 I__4832 (
            .O(N__25242),
            .I(\QuadInstance4.Quad_RNIO30S1Z0Z_9 ));
    CascadeMux I__4831 (
            .O(N__25239),
            .I(N__25236));
    InMux I__4830 (
            .O(N__25236),
            .I(N__25233));
    LocalMux I__4829 (
            .O(N__25233),
            .I(N__25230));
    Span4Mux_s2_v I__4828 (
            .O(N__25230),
            .I(N__25227));
    Odrv4 I__4827 (
            .O(N__25227),
            .I(\QuadInstance4.Quad_RNIM10S1Z0Z_7 ));
    CascadeMux I__4826 (
            .O(N__25224),
            .I(N__25221));
    InMux I__4825 (
            .O(N__25221),
            .I(N__25218));
    LocalMux I__4824 (
            .O(N__25218),
            .I(N__25215));
    Span4Mux_h I__4823 (
            .O(N__25215),
            .I(N__25211));
    InMux I__4822 (
            .O(N__25214),
            .I(N__25208));
    Span4Mux_h I__4821 (
            .O(N__25211),
            .I(N__25205));
    LocalMux I__4820 (
            .O(N__25208),
            .I(N__25202));
    Odrv4 I__4819 (
            .O(N__25205),
            .I(dataRead4_15));
    Odrv4 I__4818 (
            .O(N__25202),
            .I(dataRead4_15));
    InMux I__4817 (
            .O(N__25197),
            .I(N__25194));
    LocalMux I__4816 (
            .O(N__25194),
            .I(N__25191));
    Odrv4 I__4815 (
            .O(N__25191),
            .I(OutReg_0_5_i_m3_ns_1_15));
    InMux I__4814 (
            .O(N__25188),
            .I(\QuadInstance4.un1_Quad_cry_13 ));
    InMux I__4813 (
            .O(N__25185),
            .I(N__25182));
    LocalMux I__4812 (
            .O(N__25182),
            .I(N__25179));
    Span4Mux_v I__4811 (
            .O(N__25179),
            .I(N__25176));
    Span4Mux_h I__4810 (
            .O(N__25176),
            .I(N__25173));
    Odrv4 I__4809 (
            .O(N__25173),
            .I(\QuadInstance4.un1_Quad_axb_15 ));
    InMux I__4808 (
            .O(N__25170),
            .I(\QuadInstance4.un1_Quad_cry_14 ));
    InMux I__4807 (
            .O(N__25167),
            .I(N__25164));
    LocalMux I__4806 (
            .O(N__25164),
            .I(N__25161));
    Odrv4 I__4805 (
            .O(N__25161),
            .I(\QuadInstance4.Quad_RNO_0_4_6 ));
    CascadeMux I__4804 (
            .O(N__25158),
            .I(N__25155));
    InMux I__4803 (
            .O(N__25155),
            .I(N__25152));
    LocalMux I__4802 (
            .O(N__25152),
            .I(N__25149));
    Odrv4 I__4801 (
            .O(N__25149),
            .I(\QuadInstance4.Quad_RNIL00S1Z0Z_6 ));
    CascadeMux I__4800 (
            .O(N__25146),
            .I(N__25143));
    InMux I__4799 (
            .O(N__25143),
            .I(N__25140));
    LocalMux I__4798 (
            .O(N__25140),
            .I(\QuadInstance4.Quad_RNI06TL1Z0Z_10 ));
    CascadeMux I__4797 (
            .O(N__25137),
            .I(N__25134));
    InMux I__4796 (
            .O(N__25134),
            .I(N__25131));
    LocalMux I__4795 (
            .O(N__25131),
            .I(\QuadInstance4.Quad_RNI17TL1Z0Z_11 ));
    InMux I__4794 (
            .O(N__25128),
            .I(N__25125));
    LocalMux I__4793 (
            .O(N__25125),
            .I(\QuadInstance4.Quad_RNO_0_4_11 ));
    CascadeMux I__4792 (
            .O(N__25122),
            .I(N__25119));
    InMux I__4791 (
            .O(N__25119),
            .I(N__25116));
    LocalMux I__4790 (
            .O(N__25116),
            .I(N__25112));
    CascadeMux I__4789 (
            .O(N__25115),
            .I(N__25109));
    Span4Mux_v I__4788 (
            .O(N__25112),
            .I(N__25105));
    InMux I__4787 (
            .O(N__25109),
            .I(N__25102));
    InMux I__4786 (
            .O(N__25108),
            .I(N__25099));
    Span4Mux_h I__4785 (
            .O(N__25105),
            .I(N__25096));
    LocalMux I__4784 (
            .O(N__25102),
            .I(dataRead4_11));
    LocalMux I__4783 (
            .O(N__25099),
            .I(dataRead4_11));
    Odrv4 I__4782 (
            .O(N__25096),
            .I(dataRead4_11));
    CascadeMux I__4781 (
            .O(N__25089),
            .I(N__25084));
    CascadeMux I__4780 (
            .O(N__25088),
            .I(N__25081));
    InMux I__4779 (
            .O(N__25087),
            .I(N__25078));
    InMux I__4778 (
            .O(N__25084),
            .I(N__25075));
    InMux I__4777 (
            .O(N__25081),
            .I(N__25072));
    LocalMux I__4776 (
            .O(N__25078),
            .I(N__25069));
    LocalMux I__4775 (
            .O(N__25075),
            .I(dataRead4_6));
    LocalMux I__4774 (
            .O(N__25072),
            .I(dataRead4_6));
    Odrv4 I__4773 (
            .O(N__25069),
            .I(dataRead4_6));
    InMux I__4772 (
            .O(N__25062),
            .I(\QuadInstance4.un1_Quad_cry_4 ));
    InMux I__4771 (
            .O(N__25059),
            .I(\QuadInstance4.un1_Quad_cry_5 ));
    InMux I__4770 (
            .O(N__25056),
            .I(\QuadInstance4.un1_Quad_cry_6 ));
    InMux I__4769 (
            .O(N__25053),
            .I(bfn_15_4_0_));
    InMux I__4768 (
            .O(N__25050),
            .I(N__25047));
    LocalMux I__4767 (
            .O(N__25047),
            .I(N__25044));
    Span4Mux_v I__4766 (
            .O(N__25044),
            .I(N__25041));
    Span4Mux_h I__4765 (
            .O(N__25041),
            .I(N__25038));
    Odrv4 I__4764 (
            .O(N__25038),
            .I(\QuadInstance4.Quad_RNO_0_4_9 ));
    InMux I__4763 (
            .O(N__25035),
            .I(\QuadInstance4.un1_Quad_cry_8 ));
    InMux I__4762 (
            .O(N__25032),
            .I(\QuadInstance4.un1_Quad_cry_9 ));
    InMux I__4761 (
            .O(N__25029),
            .I(\QuadInstance4.un1_Quad_cry_10 ));
    InMux I__4760 (
            .O(N__25026),
            .I(\QuadInstance4.un1_Quad_cry_11 ));
    InMux I__4759 (
            .O(N__25023),
            .I(\QuadInstance4.un1_Quad_cry_12 ));
    InMux I__4758 (
            .O(N__25020),
            .I(N__25017));
    LocalMux I__4757 (
            .O(N__25017),
            .I(N__25014));
    Span4Mux_s3_v I__4756 (
            .O(N__25014),
            .I(N__25011));
    Span4Mux_v I__4755 (
            .O(N__25011),
            .I(N__25008));
    Span4Mux_v I__4754 (
            .O(N__25008),
            .I(N__25005));
    Odrv4 I__4753 (
            .O(N__25005),
            .I(\PWMInstance4.un1_PWMPulseWidthCount_0_I_39_c_RNO_3 ));
    InMux I__4752 (
            .O(N__25002),
            .I(N__24999));
    LocalMux I__4751 (
            .O(N__24999),
            .I(N__24996));
    Span4Mux_h I__4750 (
            .O(N__24996),
            .I(N__24993));
    Sp12to4 I__4749 (
            .O(N__24993),
            .I(N__24990));
    Span12Mux_s6_v I__4748 (
            .O(N__24990),
            .I(N__24987));
    Odrv12 I__4747 (
            .O(N__24987),
            .I(\PWMInstance4.un1_PWMPulseWidthCount_0_I_21_c_RNO_3 ));
    InMux I__4746 (
            .O(N__24984),
            .I(bfn_15_2_0_));
    IoInMux I__4745 (
            .O(N__24981),
            .I(N__24978));
    LocalMux I__4744 (
            .O(N__24978),
            .I(N__24975));
    IoSpan4Mux I__4743 (
            .O(N__24975),
            .I(N__24972));
    Span4Mux_s2_v I__4742 (
            .O(N__24972),
            .I(N__24969));
    Span4Mux_v I__4741 (
            .O(N__24969),
            .I(N__24966));
    Sp12to4 I__4740 (
            .O(N__24966),
            .I(N__24963));
    Span12Mux_v I__4739 (
            .O(N__24963),
            .I(N__24959));
    InMux I__4738 (
            .O(N__24962),
            .I(N__24956));
    Odrv12 I__4737 (
            .O(N__24959),
            .I(PWM4_c));
    LocalMux I__4736 (
            .O(N__24956),
            .I(PWM4_c));
    InMux I__4735 (
            .O(N__24951),
            .I(N__24948));
    LocalMux I__4734 (
            .O(N__24948),
            .I(N__24945));
    Span4Mux_h I__4733 (
            .O(N__24945),
            .I(N__24942));
    Odrv4 I__4732 (
            .O(N__24942),
            .I(\QuadInstance4.Quad_RNO_0_3_1 ));
    InMux I__4731 (
            .O(N__24939),
            .I(\QuadInstance4.un1_Quad_cry_0 ));
    InMux I__4730 (
            .O(N__24936),
            .I(\QuadInstance4.un1_Quad_cry_1 ));
    InMux I__4729 (
            .O(N__24933),
            .I(\QuadInstance4.un1_Quad_cry_2 ));
    InMux I__4728 (
            .O(N__24930),
            .I(N__24927));
    LocalMux I__4727 (
            .O(N__24927),
            .I(N__24924));
    Span4Mux_h I__4726 (
            .O(N__24924),
            .I(N__24921));
    Odrv4 I__4725 (
            .O(N__24921),
            .I(\QuadInstance4.Quad_RNO_0_4_4 ));
    InMux I__4724 (
            .O(N__24918),
            .I(\QuadInstance4.un1_Quad_cry_3 ));
    InMux I__4723 (
            .O(N__24915),
            .I(N__24911));
    InMux I__4722 (
            .O(N__24914),
            .I(N__24907));
    LocalMux I__4721 (
            .O(N__24911),
            .I(N__24904));
    InMux I__4720 (
            .O(N__24910),
            .I(N__24901));
    LocalMux I__4719 (
            .O(N__24907),
            .I(\PWMInstance4.periodCounterZ0Z_14 ));
    Odrv4 I__4718 (
            .O(N__24904),
            .I(\PWMInstance4.periodCounterZ0Z_14 ));
    LocalMux I__4717 (
            .O(N__24901),
            .I(\PWMInstance4.periodCounterZ0Z_14 ));
    InMux I__4716 (
            .O(N__24894),
            .I(\PWMInstance4.un1_periodCounter_2_cry_13 ));
    InMux I__4715 (
            .O(N__24891),
            .I(\PWMInstance4.un1_periodCounter_2_cry_14 ));
    InMux I__4714 (
            .O(N__24888),
            .I(bfn_14_18_0_));
    InMux I__4713 (
            .O(N__24885),
            .I(N__24882));
    LocalMux I__4712 (
            .O(N__24882),
            .I(N__24879));
    Span4Mux_s2_v I__4711 (
            .O(N__24879),
            .I(N__24876));
    Span4Mux_v I__4710 (
            .O(N__24876),
            .I(N__24873));
    Span4Mux_v I__4709 (
            .O(N__24873),
            .I(N__24870));
    Odrv4 I__4708 (
            .O(N__24870),
            .I(\PWMInstance4.un1_PWMPulseWidthCount_0_I_9_c_RNO_3 ));
    InMux I__4707 (
            .O(N__24867),
            .I(N__24864));
    LocalMux I__4706 (
            .O(N__24864),
            .I(N__24861));
    Span12Mux_h I__4705 (
            .O(N__24861),
            .I(N__24858));
    Span12Mux_v I__4704 (
            .O(N__24858),
            .I(N__24855));
    Odrv12 I__4703 (
            .O(N__24855),
            .I(\PWMInstance4.un1_PWMPulseWidthCount_0_I_15_c_RNO_3 ));
    InMux I__4702 (
            .O(N__24852),
            .I(N__24849));
    LocalMux I__4701 (
            .O(N__24849),
            .I(N__24846));
    Span4Mux_h I__4700 (
            .O(N__24846),
            .I(N__24843));
    Sp12to4 I__4699 (
            .O(N__24843),
            .I(N__24840));
    Span12Mux_s9_v I__4698 (
            .O(N__24840),
            .I(N__24837));
    Odrv12 I__4697 (
            .O(N__24837),
            .I(\PWMInstance4.un1_PWMPulseWidthCount_0_I_33_c_RNO_3 ));
    CascadeMux I__4696 (
            .O(N__24834),
            .I(N__24829));
    InMux I__4695 (
            .O(N__24833),
            .I(N__24826));
    InMux I__4694 (
            .O(N__24832),
            .I(N__24823));
    InMux I__4693 (
            .O(N__24829),
            .I(N__24820));
    LocalMux I__4692 (
            .O(N__24826),
            .I(\PWMInstance4.periodCounterZ0Z_5 ));
    LocalMux I__4691 (
            .O(N__24823),
            .I(\PWMInstance4.periodCounterZ0Z_5 ));
    LocalMux I__4690 (
            .O(N__24820),
            .I(\PWMInstance4.periodCounterZ0Z_5 ));
    InMux I__4689 (
            .O(N__24813),
            .I(\PWMInstance4.un1_periodCounter_2_cry_4 ));
    InMux I__4688 (
            .O(N__24810),
            .I(\PWMInstance4.un1_periodCounter_2_cry_5 ));
    InMux I__4687 (
            .O(N__24807),
            .I(\PWMInstance4.un1_periodCounter_2_cry_6 ));
    InMux I__4686 (
            .O(N__24804),
            .I(bfn_14_17_0_));
    InMux I__4685 (
            .O(N__24801),
            .I(\PWMInstance4.un1_periodCounter_2_cry_8 ));
    InMux I__4684 (
            .O(N__24798),
            .I(N__24793));
    InMux I__4683 (
            .O(N__24797),
            .I(N__24788));
    InMux I__4682 (
            .O(N__24796),
            .I(N__24788));
    LocalMux I__4681 (
            .O(N__24793),
            .I(\PWMInstance4.periodCounterZ0Z_10 ));
    LocalMux I__4680 (
            .O(N__24788),
            .I(\PWMInstance4.periodCounterZ0Z_10 ));
    InMux I__4679 (
            .O(N__24783),
            .I(\PWMInstance4.un1_periodCounter_2_cry_9 ));
    CascadeMux I__4678 (
            .O(N__24780),
            .I(N__24777));
    InMux I__4677 (
            .O(N__24777),
            .I(N__24772));
    CascadeMux I__4676 (
            .O(N__24776),
            .I(N__24769));
    InMux I__4675 (
            .O(N__24775),
            .I(N__24766));
    LocalMux I__4674 (
            .O(N__24772),
            .I(N__24763));
    InMux I__4673 (
            .O(N__24769),
            .I(N__24760));
    LocalMux I__4672 (
            .O(N__24766),
            .I(\PWMInstance4.periodCounterZ0Z_11 ));
    Odrv4 I__4671 (
            .O(N__24763),
            .I(\PWMInstance4.periodCounterZ0Z_11 ));
    LocalMux I__4670 (
            .O(N__24760),
            .I(\PWMInstance4.periodCounterZ0Z_11 ));
    InMux I__4669 (
            .O(N__24753),
            .I(\PWMInstance4.un1_periodCounter_2_cry_10 ));
    InMux I__4668 (
            .O(N__24750),
            .I(N__24746));
    InMux I__4667 (
            .O(N__24749),
            .I(N__24742));
    LocalMux I__4666 (
            .O(N__24746),
            .I(N__24739));
    InMux I__4665 (
            .O(N__24745),
            .I(N__24736));
    LocalMux I__4664 (
            .O(N__24742),
            .I(\PWMInstance4.periodCounterZ0Z_12 ));
    Odrv4 I__4663 (
            .O(N__24739),
            .I(\PWMInstance4.periodCounterZ0Z_12 ));
    LocalMux I__4662 (
            .O(N__24736),
            .I(\PWMInstance4.periodCounterZ0Z_12 ));
    InMux I__4661 (
            .O(N__24729),
            .I(\PWMInstance4.un1_periodCounter_2_cry_11 ));
    InMux I__4660 (
            .O(N__24726),
            .I(\PWMInstance4.un1_periodCounter_2_cry_12 ));
    InMux I__4659 (
            .O(N__24723),
            .I(N__24720));
    LocalMux I__4658 (
            .O(N__24720),
            .I(\PWMInstance4.PWMPulseWidthCountZ0Z_14 ));
    InMux I__4657 (
            .O(N__24717),
            .I(N__24714));
    LocalMux I__4656 (
            .O(N__24714),
            .I(\PWMInstance4.PWMPulseWidthCountZ0Z_15 ));
    InMux I__4655 (
            .O(N__24711),
            .I(N__24708));
    LocalMux I__4654 (
            .O(N__24708),
            .I(\PWMInstance4.PWMPulseWidthCountZ0Z_12 ));
    InMux I__4653 (
            .O(N__24705),
            .I(N__24702));
    LocalMux I__4652 (
            .O(N__24702),
            .I(\PWMInstance4.PWMPulseWidthCountZ0Z_13 ));
    InMux I__4651 (
            .O(N__24699),
            .I(\PWMInstance4.un1_periodCounter_2_cry_0 ));
    InMux I__4650 (
            .O(N__24696),
            .I(N__24691));
    InMux I__4649 (
            .O(N__24695),
            .I(N__24688));
    InMux I__4648 (
            .O(N__24694),
            .I(N__24685));
    LocalMux I__4647 (
            .O(N__24691),
            .I(\PWMInstance4.periodCounterZ0Z_2 ));
    LocalMux I__4646 (
            .O(N__24688),
            .I(\PWMInstance4.periodCounterZ0Z_2 ));
    LocalMux I__4645 (
            .O(N__24685),
            .I(\PWMInstance4.periodCounterZ0Z_2 ));
    InMux I__4644 (
            .O(N__24678),
            .I(\PWMInstance4.un1_periodCounter_2_cry_1 ));
    CascadeMux I__4643 (
            .O(N__24675),
            .I(N__24670));
    InMux I__4642 (
            .O(N__24674),
            .I(N__24667));
    InMux I__4641 (
            .O(N__24673),
            .I(N__24662));
    InMux I__4640 (
            .O(N__24670),
            .I(N__24662));
    LocalMux I__4639 (
            .O(N__24667),
            .I(\PWMInstance4.periodCounterZ0Z_3 ));
    LocalMux I__4638 (
            .O(N__24662),
            .I(\PWMInstance4.periodCounterZ0Z_3 ));
    InMux I__4637 (
            .O(N__24657),
            .I(\PWMInstance4.un1_periodCounter_2_cry_2 ));
    InMux I__4636 (
            .O(N__24654),
            .I(N__24649));
    InMux I__4635 (
            .O(N__24653),
            .I(N__24644));
    InMux I__4634 (
            .O(N__24652),
            .I(N__24644));
    LocalMux I__4633 (
            .O(N__24649),
            .I(\PWMInstance4.periodCounterZ0Z_4 ));
    LocalMux I__4632 (
            .O(N__24644),
            .I(\PWMInstance4.periodCounterZ0Z_4 ));
    InMux I__4631 (
            .O(N__24639),
            .I(\PWMInstance4.un1_periodCounter_2_cry_3 ));
    InMux I__4630 (
            .O(N__24636),
            .I(N__24629));
    InMux I__4629 (
            .O(N__24635),
            .I(N__24629));
    InMux I__4628 (
            .O(N__24634),
            .I(N__24626));
    LocalMux I__4627 (
            .O(N__24629),
            .I(pwmWriteZ0Z_3));
    LocalMux I__4626 (
            .O(N__24626),
            .I(pwmWriteZ0Z_3));
    InMux I__4625 (
            .O(N__24621),
            .I(N__24615));
    InMux I__4624 (
            .O(N__24620),
            .I(N__24615));
    LocalMux I__4623 (
            .O(N__24615),
            .I(pwmWrite_fastZ0Z_3));
    CascadeMux I__4622 (
            .O(N__24612),
            .I(N__24608));
    CascadeMux I__4621 (
            .O(N__24611),
            .I(N__24605));
    InMux I__4620 (
            .O(N__24608),
            .I(N__24594));
    InMux I__4619 (
            .O(N__24605),
            .I(N__24594));
    InMux I__4618 (
            .O(N__24604),
            .I(N__24594));
    InMux I__4617 (
            .O(N__24603),
            .I(N__24594));
    LocalMux I__4616 (
            .O(N__24594),
            .I(\PWMInstance3.clkCountZ0Z_1 ));
    InMux I__4615 (
            .O(N__24591),
            .I(N__24579));
    InMux I__4614 (
            .O(N__24590),
            .I(N__24579));
    InMux I__4613 (
            .O(N__24589),
            .I(N__24579));
    InMux I__4612 (
            .O(N__24588),
            .I(N__24579));
    LocalMux I__4611 (
            .O(N__24579),
            .I(\PWMInstance3.clkCountZ0Z_0 ));
    CascadeMux I__4610 (
            .O(N__24576),
            .I(\PWMInstance3.un1_periodCounter12_1_0_a2_0_6_cascade_ ));
    CascadeMux I__4609 (
            .O(N__24573),
            .I(\PWMInstance3.un1_periodCounter12_1_0_a2_0_14_cascade_ ));
    InMux I__4608 (
            .O(N__24570),
            .I(N__24567));
    LocalMux I__4607 (
            .O(N__24567),
            .I(N__24564));
    Span4Mux_v I__4606 (
            .O(N__24564),
            .I(N__24561));
    Odrv4 I__4605 (
            .O(N__24561),
            .I(\PWMInstance6.PWMPulseWidthCountZ0Z_9 ));
    CEMux I__4604 (
            .O(N__24558),
            .I(N__24553));
    CEMux I__4603 (
            .O(N__24557),
            .I(N__24549));
    CEMux I__4602 (
            .O(N__24556),
            .I(N__24546));
    LocalMux I__4601 (
            .O(N__24553),
            .I(N__24543));
    CEMux I__4600 (
            .O(N__24552),
            .I(N__24540));
    LocalMux I__4599 (
            .O(N__24549),
            .I(N__24536));
    LocalMux I__4598 (
            .O(N__24546),
            .I(N__24533));
    Span4Mux_v I__4597 (
            .O(N__24543),
            .I(N__24530));
    LocalMux I__4596 (
            .O(N__24540),
            .I(N__24527));
    CEMux I__4595 (
            .O(N__24539),
            .I(N__24524));
    Span4Mux_v I__4594 (
            .O(N__24536),
            .I(N__24521));
    Span4Mux_h I__4593 (
            .O(N__24533),
            .I(N__24518));
    Span4Mux_h I__4592 (
            .O(N__24530),
            .I(N__24513));
    Span4Mux_h I__4591 (
            .O(N__24527),
            .I(N__24513));
    LocalMux I__4590 (
            .O(N__24524),
            .I(N__24510));
    Span4Mux_h I__4589 (
            .O(N__24521),
            .I(N__24507));
    Odrv4 I__4588 (
            .O(N__24518),
            .I(\PWMInstance6.pwmWrite_0_6 ));
    Odrv4 I__4587 (
            .O(N__24513),
            .I(\PWMInstance6.pwmWrite_0_6 ));
    Odrv12 I__4586 (
            .O(N__24510),
            .I(\PWMInstance6.pwmWrite_0_6 ));
    Odrv4 I__4585 (
            .O(N__24507),
            .I(\PWMInstance6.pwmWrite_0_6 ));
    InMux I__4584 (
            .O(N__24498),
            .I(N__24495));
    LocalMux I__4583 (
            .O(N__24495),
            .I(\PWMInstance4.PWMPulseWidthCountZ0Z_3 ));
    InMux I__4582 (
            .O(N__24492),
            .I(N__24489));
    LocalMux I__4581 (
            .O(N__24489),
            .I(\PWMInstance4.PWMPulseWidthCountZ0Z_2 ));
    InMux I__4580 (
            .O(N__24486),
            .I(N__24482));
    InMux I__4579 (
            .O(N__24485),
            .I(N__24479));
    LocalMux I__4578 (
            .O(N__24482),
            .I(data_receivedZ0Z_8));
    LocalMux I__4577 (
            .O(N__24479),
            .I(data_receivedZ0Z_8));
    InMux I__4576 (
            .O(N__24474),
            .I(N__24470));
    InMux I__4575 (
            .O(N__24473),
            .I(N__24467));
    LocalMux I__4574 (
            .O(N__24470),
            .I(data_receivedZ0Z_9));
    LocalMux I__4573 (
            .O(N__24467),
            .I(data_receivedZ0Z_9));
    CEMux I__4572 (
            .O(N__24462),
            .I(N__24458));
    CEMux I__4571 (
            .O(N__24461),
            .I(N__24455));
    LocalMux I__4570 (
            .O(N__24458),
            .I(N_870_i));
    LocalMux I__4569 (
            .O(N__24455),
            .I(N_870_i));
    InMux I__4568 (
            .O(N__24450),
            .I(N__24446));
    InMux I__4567 (
            .O(N__24449),
            .I(N__24443));
    LocalMux I__4566 (
            .O(N__24446),
            .I(data_receivedZ0Z_5));
    LocalMux I__4565 (
            .O(N__24443),
            .I(data_receivedZ0Z_5));
    InMux I__4564 (
            .O(N__24438),
            .I(N__24434));
    InMux I__4563 (
            .O(N__24437),
            .I(N__24431));
    LocalMux I__4562 (
            .O(N__24434),
            .I(data_receivedZ0Z_6));
    LocalMux I__4561 (
            .O(N__24431),
            .I(data_receivedZ0Z_6));
    InMux I__4560 (
            .O(N__24426),
            .I(N__24422));
    InMux I__4559 (
            .O(N__24425),
            .I(N__24419));
    LocalMux I__4558 (
            .O(N__24422),
            .I(data_receivedZ0Z_7));
    LocalMux I__4557 (
            .O(N__24419),
            .I(data_receivedZ0Z_7));
    InMux I__4556 (
            .O(N__24414),
            .I(N__24411));
    LocalMux I__4555 (
            .O(N__24411),
            .I(N__24407));
    InMux I__4554 (
            .O(N__24410),
            .I(N__24403));
    Span4Mux_v I__4553 (
            .O(N__24407),
            .I(N__24400));
    InMux I__4552 (
            .O(N__24406),
            .I(N__24397));
    LocalMux I__4551 (
            .O(N__24403),
            .I(N__24394));
    Span4Mux_v I__4550 (
            .O(N__24400),
            .I(N__24389));
    LocalMux I__4549 (
            .O(N__24397),
            .I(N__24389));
    Span4Mux_h I__4548 (
            .O(N__24394),
            .I(N__24386));
    Span4Mux_h I__4547 (
            .O(N__24389),
            .I(N__24383));
    Span4Mux_v I__4546 (
            .O(N__24386),
            .I(N__24380));
    Odrv4 I__4545 (
            .O(N__24383),
            .I(dataRead2_3));
    Odrv4 I__4544 (
            .O(N__24380),
            .I(dataRead2_3));
    InMux I__4543 (
            .O(N__24375),
            .I(N__24371));
    CascadeMux I__4542 (
            .O(N__24374),
            .I(N__24368));
    LocalMux I__4541 (
            .O(N__24371),
            .I(N__24364));
    InMux I__4540 (
            .O(N__24368),
            .I(N__24361));
    InMux I__4539 (
            .O(N__24367),
            .I(N__24358));
    Span4Mux_h I__4538 (
            .O(N__24364),
            .I(N__24355));
    LocalMux I__4537 (
            .O(N__24361),
            .I(N__24352));
    LocalMux I__4536 (
            .O(N__24358),
            .I(N__24349));
    Span4Mux_v I__4535 (
            .O(N__24355),
            .I(N__24346));
    Span4Mux_h I__4534 (
            .O(N__24352),
            .I(N__24341));
    Span4Mux_h I__4533 (
            .O(N__24349),
            .I(N__24341));
    Odrv4 I__4532 (
            .O(N__24346),
            .I(dataRead3_3));
    Odrv4 I__4531 (
            .O(N__24341),
            .I(dataRead3_3));
    InMux I__4530 (
            .O(N__24336),
            .I(N__24332));
    InMux I__4529 (
            .O(N__24335),
            .I(N__24329));
    LocalMux I__4528 (
            .O(N__24332),
            .I(N__24326));
    LocalMux I__4527 (
            .O(N__24329),
            .I(N__24323));
    Span4Mux_h I__4526 (
            .O(N__24326),
            .I(N__24320));
    Odrv4 I__4525 (
            .O(N__24323),
            .I(dataRead3_15));
    Odrv4 I__4524 (
            .O(N__24320),
            .I(dataRead3_15));
    InMux I__4523 (
            .O(N__24315),
            .I(N__24311));
    CascadeMux I__4522 (
            .O(N__24314),
            .I(N__24308));
    LocalMux I__4521 (
            .O(N__24311),
            .I(N__24305));
    InMux I__4520 (
            .O(N__24308),
            .I(N__24302));
    Span4Mux_h I__4519 (
            .O(N__24305),
            .I(N__24299));
    LocalMux I__4518 (
            .O(N__24302),
            .I(N__24294));
    Span4Mux_h I__4517 (
            .O(N__24299),
            .I(N__24294));
    Odrv4 I__4516 (
            .O(N__24294),
            .I(dataRead2_15));
    InMux I__4515 (
            .O(N__24291),
            .I(N__24287));
    InMux I__4514 (
            .O(N__24290),
            .I(N__24284));
    LocalMux I__4513 (
            .O(N__24287),
            .I(N__24281));
    LocalMux I__4512 (
            .O(N__24284),
            .I(N__24276));
    Span4Mux_h I__4511 (
            .O(N__24281),
            .I(N__24276));
    Odrv4 I__4510 (
            .O(N__24276),
            .I(dataRead7_15));
    CascadeMux I__4509 (
            .O(N__24273),
            .I(N__24270));
    InMux I__4508 (
            .O(N__24270),
            .I(N__24266));
    InMux I__4507 (
            .O(N__24269),
            .I(N__24263));
    LocalMux I__4506 (
            .O(N__24266),
            .I(N__24260));
    LocalMux I__4505 (
            .O(N__24263),
            .I(N__24257));
    Span4Mux_v I__4504 (
            .O(N__24260),
            .I(N__24252));
    Span4Mux_h I__4503 (
            .O(N__24257),
            .I(N__24252));
    Odrv4 I__4502 (
            .O(N__24252),
            .I(dataRead6_15));
    CascadeMux I__4501 (
            .O(N__24249),
            .I(OutReg_0_4_i_m3_ns_1_15_cascade_));
    InMux I__4500 (
            .O(N__24246),
            .I(N__24243));
    LocalMux I__4499 (
            .O(N__24243),
            .I(N__24239));
    InMux I__4498 (
            .O(N__24242),
            .I(N__24236));
    Span4Mux_h I__4497 (
            .O(N__24239),
            .I(N__24233));
    LocalMux I__4496 (
            .O(N__24236),
            .I(dataRead5_15));
    Odrv4 I__4495 (
            .O(N__24233),
            .I(dataRead5_15));
    CascadeMux I__4494 (
            .O(N__24228),
            .I(N__24224));
    InMux I__4493 (
            .O(N__24227),
            .I(N__24221));
    InMux I__4492 (
            .O(N__24224),
            .I(N__24218));
    LocalMux I__4491 (
            .O(N__24221),
            .I(N__24213));
    LocalMux I__4490 (
            .O(N__24218),
            .I(N__24213));
    Odrv4 I__4489 (
            .O(N__24213),
            .I(dataRead1_15));
    CascadeMux I__4488 (
            .O(N__24210),
            .I(N__24205));
    CascadeMux I__4487 (
            .O(N__24209),
            .I(N__24202));
    InMux I__4486 (
            .O(N__24208),
            .I(N__24183));
    InMux I__4485 (
            .O(N__24205),
            .I(N__24183));
    InMux I__4484 (
            .O(N__24202),
            .I(N__24183));
    InMux I__4483 (
            .O(N__24201),
            .I(N__24183));
    InMux I__4482 (
            .O(N__24200),
            .I(N__24183));
    InMux I__4481 (
            .O(N__24199),
            .I(N__24183));
    CascadeMux I__4480 (
            .O(N__24198),
            .I(N__24175));
    CascadeMux I__4479 (
            .O(N__24197),
            .I(N__24170));
    InMux I__4478 (
            .O(N__24196),
            .I(N__24167));
    LocalMux I__4477 (
            .O(N__24183),
            .I(N__24164));
    InMux I__4476 (
            .O(N__24182),
            .I(N__24157));
    InMux I__4475 (
            .O(N__24181),
            .I(N__24157));
    InMux I__4474 (
            .O(N__24180),
            .I(N__24157));
    InMux I__4473 (
            .O(N__24179),
            .I(N__24144));
    InMux I__4472 (
            .O(N__24178),
            .I(N__24144));
    InMux I__4471 (
            .O(N__24175),
            .I(N__24144));
    InMux I__4470 (
            .O(N__24174),
            .I(N__24144));
    InMux I__4469 (
            .O(N__24173),
            .I(N__24144));
    InMux I__4468 (
            .O(N__24170),
            .I(N__24144));
    LocalMux I__4467 (
            .O(N__24167),
            .I(\QuadInstance1.count_enable ));
    Odrv4 I__4466 (
            .O(N__24164),
            .I(\QuadInstance1.count_enable ));
    LocalMux I__4465 (
            .O(N__24157),
            .I(\QuadInstance1.count_enable ));
    LocalMux I__4464 (
            .O(N__24144),
            .I(\QuadInstance1.count_enable ));
    InMux I__4463 (
            .O(N__24135),
            .I(N__24132));
    LocalMux I__4462 (
            .O(N__24132),
            .I(\QuadInstance1.Quad_RNO_0_1_12 ));
    InMux I__4461 (
            .O(N__24129),
            .I(N__24125));
    CascadeMux I__4460 (
            .O(N__24128),
            .I(N__24122));
    LocalMux I__4459 (
            .O(N__24125),
            .I(N__24118));
    InMux I__4458 (
            .O(N__24122),
            .I(N__24115));
    InMux I__4457 (
            .O(N__24121),
            .I(N__24112));
    Span4Mux_v I__4456 (
            .O(N__24118),
            .I(N__24109));
    LocalMux I__4455 (
            .O(N__24115),
            .I(dataRead1_12));
    LocalMux I__4454 (
            .O(N__24112),
            .I(dataRead1_12));
    Odrv4 I__4453 (
            .O(N__24109),
            .I(dataRead1_12));
    InMux I__4452 (
            .O(N__24102),
            .I(N__24092));
    InMux I__4451 (
            .O(N__24101),
            .I(N__24087));
    InMux I__4450 (
            .O(N__24100),
            .I(N__24087));
    CascadeMux I__4449 (
            .O(N__24099),
            .I(N__24081));
    InMux I__4448 (
            .O(N__24098),
            .I(N__24077));
    InMux I__4447 (
            .O(N__24097),
            .I(N__24072));
    InMux I__4446 (
            .O(N__24096),
            .I(N__24072));
    InMux I__4445 (
            .O(N__24095),
            .I(N__24069));
    LocalMux I__4444 (
            .O(N__24092),
            .I(N__24066));
    LocalMux I__4443 (
            .O(N__24087),
            .I(N__24063));
    InMux I__4442 (
            .O(N__24086),
            .I(N__24060));
    CascadeMux I__4441 (
            .O(N__24085),
            .I(N__24056));
    CascadeMux I__4440 (
            .O(N__24084),
            .I(N__24053));
    InMux I__4439 (
            .O(N__24081),
            .I(N__24045));
    InMux I__4438 (
            .O(N__24080),
            .I(N__24045));
    LocalMux I__4437 (
            .O(N__24077),
            .I(N__24042));
    LocalMux I__4436 (
            .O(N__24072),
            .I(N__24037));
    LocalMux I__4435 (
            .O(N__24069),
            .I(N__24037));
    Span4Mux_v I__4434 (
            .O(N__24066),
            .I(N__24032));
    Span4Mux_v I__4433 (
            .O(N__24063),
            .I(N__24032));
    LocalMux I__4432 (
            .O(N__24060),
            .I(N__24029));
    InMux I__4431 (
            .O(N__24059),
            .I(N__24018));
    InMux I__4430 (
            .O(N__24056),
            .I(N__24011));
    InMux I__4429 (
            .O(N__24053),
            .I(N__24011));
    InMux I__4428 (
            .O(N__24052),
            .I(N__24011));
    InMux I__4427 (
            .O(N__24051),
            .I(N__24001));
    InMux I__4426 (
            .O(N__24050),
            .I(N__23998));
    LocalMux I__4425 (
            .O(N__24045),
            .I(N__23993));
    Span4Mux_v I__4424 (
            .O(N__24042),
            .I(N__23993));
    Span4Mux_h I__4423 (
            .O(N__24037),
            .I(N__23990));
    Sp12to4 I__4422 (
            .O(N__24032),
            .I(N__23985));
    Span12Mux_v I__4421 (
            .O(N__24029),
            .I(N__23985));
    InMux I__4420 (
            .O(N__24028),
            .I(N__23968));
    InMux I__4419 (
            .O(N__24027),
            .I(N__23968));
    InMux I__4418 (
            .O(N__24026),
            .I(N__23968));
    InMux I__4417 (
            .O(N__24025),
            .I(N__23968));
    InMux I__4416 (
            .O(N__24024),
            .I(N__23968));
    InMux I__4415 (
            .O(N__24023),
            .I(N__23968));
    InMux I__4414 (
            .O(N__24022),
            .I(N__23968));
    InMux I__4413 (
            .O(N__24021),
            .I(N__23968));
    LocalMux I__4412 (
            .O(N__24018),
            .I(N__23963));
    LocalMux I__4411 (
            .O(N__24011),
            .I(N__23963));
    InMux I__4410 (
            .O(N__24010),
            .I(N__23950));
    InMux I__4409 (
            .O(N__24009),
            .I(N__23950));
    InMux I__4408 (
            .O(N__24008),
            .I(N__23950));
    InMux I__4407 (
            .O(N__24007),
            .I(N__23950));
    InMux I__4406 (
            .O(N__24006),
            .I(N__23950));
    InMux I__4405 (
            .O(N__24005),
            .I(N__23950));
    InMux I__4404 (
            .O(N__24004),
            .I(N__23947));
    LocalMux I__4403 (
            .O(N__24001),
            .I(quadWriteZ0Z_1));
    LocalMux I__4402 (
            .O(N__23998),
            .I(quadWriteZ0Z_1));
    Odrv4 I__4401 (
            .O(N__23993),
            .I(quadWriteZ0Z_1));
    Odrv4 I__4400 (
            .O(N__23990),
            .I(quadWriteZ0Z_1));
    Odrv12 I__4399 (
            .O(N__23985),
            .I(quadWriteZ0Z_1));
    LocalMux I__4398 (
            .O(N__23968),
            .I(quadWriteZ0Z_1));
    Odrv4 I__4397 (
            .O(N__23963),
            .I(quadWriteZ0Z_1));
    LocalMux I__4396 (
            .O(N__23950),
            .I(quadWriteZ0Z_1));
    LocalMux I__4395 (
            .O(N__23947),
            .I(quadWriteZ0Z_1));
    InMux I__4394 (
            .O(N__23928),
            .I(N__23925));
    LocalMux I__4393 (
            .O(N__23925),
            .I(\QuadInstance1.Quad_RNO_0_1_13 ));
    InMux I__4392 (
            .O(N__23922),
            .I(N__23919));
    LocalMux I__4391 (
            .O(N__23919),
            .I(N__23914));
    InMux I__4390 (
            .O(N__23918),
            .I(N__23911));
    InMux I__4389 (
            .O(N__23917),
            .I(N__23908));
    Span4Mux_v I__4388 (
            .O(N__23914),
            .I(N__23905));
    LocalMux I__4387 (
            .O(N__23911),
            .I(dataRead1_13));
    LocalMux I__4386 (
            .O(N__23908),
            .I(dataRead1_13));
    Odrv4 I__4385 (
            .O(N__23905),
            .I(dataRead1_13));
    InMux I__4384 (
            .O(N__23898),
            .I(N__23894));
    InMux I__4383 (
            .O(N__23897),
            .I(N__23891));
    LocalMux I__4382 (
            .O(N__23894),
            .I(N__23887));
    LocalMux I__4381 (
            .O(N__23891),
            .I(N__23884));
    InMux I__4380 (
            .O(N__23890),
            .I(N__23881));
    Span4Mux_v I__4379 (
            .O(N__23887),
            .I(N__23878));
    Span4Mux_v I__4378 (
            .O(N__23884),
            .I(N__23873));
    LocalMux I__4377 (
            .O(N__23881),
            .I(N__23873));
    Odrv4 I__4376 (
            .O(N__23878),
            .I(dataRead1_1));
    Odrv4 I__4375 (
            .O(N__23873),
            .I(dataRead1_1));
    CascadeMux I__4374 (
            .O(N__23868),
            .I(N__23865));
    InMux I__4373 (
            .O(N__23865),
            .I(N__23862));
    LocalMux I__4372 (
            .O(N__23862),
            .I(N__23859));
    Span4Mux_h I__4371 (
            .O(N__23859),
            .I(N__23855));
    InMux I__4370 (
            .O(N__23858),
            .I(N__23851));
    Span4Mux_h I__4369 (
            .O(N__23855),
            .I(N__23848));
    InMux I__4368 (
            .O(N__23854),
            .I(N__23845));
    LocalMux I__4367 (
            .O(N__23851),
            .I(dataRead5_1));
    Odrv4 I__4366 (
            .O(N__23848),
            .I(dataRead5_1));
    LocalMux I__4365 (
            .O(N__23845),
            .I(dataRead5_1));
    CascadeMux I__4364 (
            .O(N__23838),
            .I(OutReg_ess_RNO_2Z0Z_1_cascade_));
    InMux I__4363 (
            .O(N__23835),
            .I(N__23831));
    InMux I__4362 (
            .O(N__23834),
            .I(N__23828));
    LocalMux I__4361 (
            .O(N__23831),
            .I(N__23822));
    LocalMux I__4360 (
            .O(N__23828),
            .I(N__23822));
    InMux I__4359 (
            .O(N__23827),
            .I(N__23819));
    Span12Mux_s7_v I__4358 (
            .O(N__23822),
            .I(N__23816));
    LocalMux I__4357 (
            .O(N__23819),
            .I(dataRead2_1));
    Odrv12 I__4356 (
            .O(N__23816),
            .I(dataRead2_1));
    InMux I__4355 (
            .O(N__23811),
            .I(N__23808));
    LocalMux I__4354 (
            .O(N__23808),
            .I(N__23804));
    InMux I__4353 (
            .O(N__23807),
            .I(N__23801));
    Span4Mux_v I__4352 (
            .O(N__23804),
            .I(N__23795));
    LocalMux I__4351 (
            .O(N__23801),
            .I(N__23795));
    InMux I__4350 (
            .O(N__23800),
            .I(N__23792));
    Odrv4 I__4349 (
            .O(N__23795),
            .I(dataRead3_1));
    LocalMux I__4348 (
            .O(N__23792),
            .I(dataRead3_1));
    InMux I__4347 (
            .O(N__23787),
            .I(N__23784));
    LocalMux I__4346 (
            .O(N__23784),
            .I(N__23779));
    InMux I__4345 (
            .O(N__23783),
            .I(N__23776));
    InMux I__4344 (
            .O(N__23782),
            .I(N__23773));
    Span4Mux_h I__4343 (
            .O(N__23779),
            .I(N__23770));
    LocalMux I__4342 (
            .O(N__23776),
            .I(N__23767));
    LocalMux I__4341 (
            .O(N__23773),
            .I(dataRead6_1));
    Odrv4 I__4340 (
            .O(N__23770),
            .I(dataRead6_1));
    Odrv4 I__4339 (
            .O(N__23767),
            .I(dataRead6_1));
    CascadeMux I__4338 (
            .O(N__23760),
            .I(OutReg_0_4_i_m3_ns_1_1_cascade_));
    InMux I__4337 (
            .O(N__23757),
            .I(N__23754));
    LocalMux I__4336 (
            .O(N__23754),
            .I(OutReg_ess_RNO_1Z0Z_1));
    InMux I__4335 (
            .O(N__23751),
            .I(N__23748));
    LocalMux I__4334 (
            .O(N__23748),
            .I(OutReg_0_5_i_m3_ns_1_1));
    InMux I__4333 (
            .O(N__23745),
            .I(N__23742));
    LocalMux I__4332 (
            .O(N__23742),
            .I(N__23738));
    InMux I__4331 (
            .O(N__23741),
            .I(N__23735));
    Span4Mux_h I__4330 (
            .O(N__23738),
            .I(N__23729));
    LocalMux I__4329 (
            .O(N__23735),
            .I(N__23729));
    InMux I__4328 (
            .O(N__23734),
            .I(N__23726));
    Span4Mux_v I__4327 (
            .O(N__23729),
            .I(N__23721));
    LocalMux I__4326 (
            .O(N__23726),
            .I(N__23721));
    Odrv4 I__4325 (
            .O(N__23721),
            .I(dataRead3_5));
    InMux I__4324 (
            .O(N__23718),
            .I(N__23714));
    InMux I__4323 (
            .O(N__23717),
            .I(N__23711));
    LocalMux I__4322 (
            .O(N__23714),
            .I(N__23707));
    LocalMux I__4321 (
            .O(N__23711),
            .I(N__23704));
    InMux I__4320 (
            .O(N__23710),
            .I(N__23701));
    Span4Mux_v I__4319 (
            .O(N__23707),
            .I(N__23696));
    Span4Mux_h I__4318 (
            .O(N__23704),
            .I(N__23696));
    LocalMux I__4317 (
            .O(N__23701),
            .I(N__23693));
    Span4Mux_h I__4316 (
            .O(N__23696),
            .I(N__23688));
    Span4Mux_h I__4315 (
            .O(N__23693),
            .I(N__23688));
    Odrv4 I__4314 (
            .O(N__23688),
            .I(dataRead2_5));
    CascadeMux I__4313 (
            .O(N__23685),
            .I(N__23682));
    InMux I__4312 (
            .O(N__23682),
            .I(N__23679));
    LocalMux I__4311 (
            .O(N__23679),
            .I(\QuadInstance1.Quad_RNIUN0OZ0Z_7 ));
    CascadeMux I__4310 (
            .O(N__23676),
            .I(N__23673));
    InMux I__4309 (
            .O(N__23673),
            .I(N__23670));
    LocalMux I__4308 (
            .O(N__23670),
            .I(\QuadInstance1.Quad_RNIPI0OZ0Z_2 ));
    CascadeMux I__4307 (
            .O(N__23667),
            .I(N__23664));
    InMux I__4306 (
            .O(N__23664),
            .I(N__23661));
    LocalMux I__4305 (
            .O(N__23661),
            .I(\QuadInstance1.Quad_RNIQJ0OZ0Z_3 ));
    CascadeMux I__4304 (
            .O(N__23658),
            .I(N__23655));
    InMux I__4303 (
            .O(N__23655),
            .I(N__23652));
    LocalMux I__4302 (
            .O(N__23652),
            .I(\QuadInstance1.Quad_RNIAR5DZ0Z_12 ));
    CascadeMux I__4301 (
            .O(N__23649),
            .I(N__23646));
    InMux I__4300 (
            .O(N__23646),
            .I(N__23643));
    LocalMux I__4299 (
            .O(N__23643),
            .I(\QuadInstance1.Quad_RNIBS5DZ0Z_13 ));
    InMux I__4298 (
            .O(N__23640),
            .I(N__23637));
    LocalMux I__4297 (
            .O(N__23637),
            .I(\QuadInstance1.Quad_RNICT5DZ0Z_14 ));
    CascadeMux I__4296 (
            .O(N__23634),
            .I(N__23631));
    InMux I__4295 (
            .O(N__23631),
            .I(N__23628));
    LocalMux I__4294 (
            .O(N__23628),
            .I(\QuadInstance1.Quad_RNIVO0OZ0Z_8 ));
    CascadeMux I__4293 (
            .O(N__23625),
            .I(N__23619));
    CascadeMux I__4292 (
            .O(N__23624),
            .I(N__23615));
    InMux I__4291 (
            .O(N__23623),
            .I(N__23599));
    InMux I__4290 (
            .O(N__23622),
            .I(N__23599));
    InMux I__4289 (
            .O(N__23619),
            .I(N__23599));
    InMux I__4288 (
            .O(N__23618),
            .I(N__23599));
    InMux I__4287 (
            .O(N__23615),
            .I(N__23599));
    CascadeMux I__4286 (
            .O(N__23614),
            .I(N__23596));
    CascadeMux I__4285 (
            .O(N__23613),
            .I(N__23592));
    CascadeMux I__4284 (
            .O(N__23612),
            .I(N__23589));
    CascadeMux I__4283 (
            .O(N__23611),
            .I(N__23585));
    CascadeMux I__4282 (
            .O(N__23610),
            .I(N__23582));
    LocalMux I__4281 (
            .O(N__23599),
            .I(N__23576));
    InMux I__4280 (
            .O(N__23596),
            .I(N__23563));
    InMux I__4279 (
            .O(N__23595),
            .I(N__23563));
    InMux I__4278 (
            .O(N__23592),
            .I(N__23563));
    InMux I__4277 (
            .O(N__23589),
            .I(N__23563));
    InMux I__4276 (
            .O(N__23588),
            .I(N__23563));
    InMux I__4275 (
            .O(N__23585),
            .I(N__23563));
    InMux I__4274 (
            .O(N__23582),
            .I(N__23554));
    InMux I__4273 (
            .O(N__23581),
            .I(N__23554));
    InMux I__4272 (
            .O(N__23580),
            .I(N__23554));
    InMux I__4271 (
            .O(N__23579),
            .I(N__23554));
    Odrv4 I__4270 (
            .O(N__23576),
            .I(\QuadInstance1.un1_count_enable_i_a2_0_1 ));
    LocalMux I__4269 (
            .O(N__23563),
            .I(\QuadInstance1.un1_count_enable_i_a2_0_1 ));
    LocalMux I__4268 (
            .O(N__23554),
            .I(\QuadInstance1.un1_count_enable_i_a2_0_1 ));
    InMux I__4267 (
            .O(N__23547),
            .I(N__23544));
    LocalMux I__4266 (
            .O(N__23544),
            .I(\QuadInstance1.un1_Quad_axb_15 ));
    CascadeMux I__4265 (
            .O(N__23541),
            .I(\QuadInstance1.count_enable_cascade_ ));
    CascadeMux I__4264 (
            .O(N__23538),
            .I(N__23535));
    InMux I__4263 (
            .O(N__23535),
            .I(N__23532));
    LocalMux I__4262 (
            .O(N__23532),
            .I(\QuadInstance1.Quad_RNIOH0OZ0Z_1 ));
    CascadeMux I__4261 (
            .O(N__23529),
            .I(N__23526));
    InMux I__4260 (
            .O(N__23526),
            .I(N__23523));
    LocalMux I__4259 (
            .O(N__23523),
            .I(\QuadInstance1.Quad_RNITM0OZ0Z_6 ));
    CascadeMux I__4258 (
            .O(N__23520),
            .I(N__23517));
    InMux I__4257 (
            .O(N__23517),
            .I(N__23514));
    LocalMux I__4256 (
            .O(N__23514),
            .I(\QuadInstance1.Quad_RNISL0OZ0Z_5 ));
    CascadeMux I__4255 (
            .O(N__23511),
            .I(N__23508));
    InMux I__4254 (
            .O(N__23508),
            .I(N__23505));
    LocalMux I__4253 (
            .O(N__23505),
            .I(\QuadInstance1.delayedCh_AZ0Z_2 ));
    InMux I__4252 (
            .O(N__23502),
            .I(N__23496));
    InMux I__4251 (
            .O(N__23501),
            .I(N__23496));
    LocalMux I__4250 (
            .O(N__23496),
            .I(\QuadInstance1.delayedCh_BZ0Z_2 ));
    InMux I__4249 (
            .O(N__23493),
            .I(N__23484));
    InMux I__4248 (
            .O(N__23492),
            .I(N__23484));
    InMux I__4247 (
            .O(N__23491),
            .I(N__23484));
    LocalMux I__4246 (
            .O(N__23484),
            .I(\QuadInstance1.delayedCh_AZ0Z_1 ));
    CascadeMux I__4245 (
            .O(N__23481),
            .I(N__23478));
    InMux I__4244 (
            .O(N__23478),
            .I(N__23475));
    LocalMux I__4243 (
            .O(N__23475),
            .I(\QuadInstance1.Quad_RNI0Q0OZ0Z_9 ));
    CascadeMux I__4242 (
            .O(N__23472),
            .I(N__23469));
    InMux I__4241 (
            .O(N__23469),
            .I(N__23466));
    LocalMux I__4240 (
            .O(N__23466),
            .I(\QuadInstance1.Quad_RNI8P5DZ0Z_10 ));
    InMux I__4239 (
            .O(N__23463),
            .I(N__23460));
    LocalMux I__4238 (
            .O(N__23460),
            .I(N__23455));
    InMux I__4237 (
            .O(N__23459),
            .I(N__23452));
    InMux I__4236 (
            .O(N__23458),
            .I(N__23445));
    Span4Mux_v I__4235 (
            .O(N__23455),
            .I(N__23441));
    LocalMux I__4234 (
            .O(N__23452),
            .I(N__23438));
    InMux I__4233 (
            .O(N__23451),
            .I(N__23435));
    InMux I__4232 (
            .O(N__23450),
            .I(N__23430));
    InMux I__4231 (
            .O(N__23449),
            .I(N__23430));
    InMux I__4230 (
            .O(N__23448),
            .I(N__23425));
    LocalMux I__4229 (
            .O(N__23445),
            .I(N__23422));
    InMux I__4228 (
            .O(N__23444),
            .I(N__23419));
    Span4Mux_h I__4227 (
            .O(N__23441),
            .I(N__23410));
    Span4Mux_v I__4226 (
            .O(N__23438),
            .I(N__23410));
    LocalMux I__4225 (
            .O(N__23435),
            .I(N__23410));
    LocalMux I__4224 (
            .O(N__23430),
            .I(N__23410));
    InMux I__4223 (
            .O(N__23429),
            .I(N__23405));
    InMux I__4222 (
            .O(N__23428),
            .I(N__23405));
    LocalMux I__4221 (
            .O(N__23425),
            .I(N__23402));
    Span4Mux_h I__4220 (
            .O(N__23422),
            .I(N__23397));
    LocalMux I__4219 (
            .O(N__23419),
            .I(N__23397));
    Span4Mux_v I__4218 (
            .O(N__23410),
            .I(N__23392));
    LocalMux I__4217 (
            .O(N__23405),
            .I(N__23392));
    Span4Mux_v I__4216 (
            .O(N__23402),
            .I(N__23388));
    Span4Mux_v I__4215 (
            .O(N__23397),
            .I(N__23385));
    Span4Mux_h I__4214 (
            .O(N__23392),
            .I(N__23382));
    InMux I__4213 (
            .O(N__23391),
            .I(N__23379));
    Odrv4 I__4212 (
            .O(N__23388),
            .I(data_received_esr_RNIMIH31Z0Z_19));
    Odrv4 I__4211 (
            .O(N__23385),
            .I(data_received_esr_RNIMIH31Z0Z_19));
    Odrv4 I__4210 (
            .O(N__23382),
            .I(data_received_esr_RNIMIH31Z0Z_19));
    LocalMux I__4209 (
            .O(N__23379),
            .I(data_received_esr_RNIMIH31Z0Z_19));
    InMux I__4208 (
            .O(N__23370),
            .I(N__23367));
    LocalMux I__4207 (
            .O(N__23367),
            .I(N__23363));
    InMux I__4206 (
            .O(N__23366),
            .I(N__23359));
    Span4Mux_v I__4205 (
            .O(N__23363),
            .I(N__23356));
    InMux I__4204 (
            .O(N__23362),
            .I(N__23353));
    LocalMux I__4203 (
            .O(N__23359),
            .I(N__23350));
    Span4Mux_v I__4202 (
            .O(N__23356),
            .I(N__23345));
    LocalMux I__4201 (
            .O(N__23353),
            .I(N__23345));
    Odrv12 I__4200 (
            .O(N__23350),
            .I(dataRead1_11));
    Odrv4 I__4199 (
            .O(N__23345),
            .I(dataRead1_11));
    CascadeMux I__4198 (
            .O(N__23340),
            .I(N__23337));
    InMux I__4197 (
            .O(N__23337),
            .I(N__23334));
    LocalMux I__4196 (
            .O(N__23334),
            .I(\QuadInstance1.Quad_RNI9Q5DZ0Z_11 ));
    InMux I__4195 (
            .O(N__23331),
            .I(N__23328));
    LocalMux I__4194 (
            .O(N__23328),
            .I(\PWMInstance4.PWMPulseWidthCountZ0Z_11 ));
    InMux I__4193 (
            .O(N__23325),
            .I(N__23322));
    LocalMux I__4192 (
            .O(N__23322),
            .I(N__23319));
    Span4Mux_h I__4191 (
            .O(N__23319),
            .I(N__23316));
    Odrv4 I__4190 (
            .O(N__23316),
            .I(ch2_B_c));
    InMux I__4189 (
            .O(N__23313),
            .I(N__23310));
    LocalMux I__4188 (
            .O(N__23310),
            .I(N__23307));
    Span4Mux_h I__4187 (
            .O(N__23307),
            .I(N__23304));
    Sp12to4 I__4186 (
            .O(N__23304),
            .I(N__23301));
    Span12Mux_v I__4185 (
            .O(N__23301),
            .I(N__23298));
    Odrv12 I__4184 (
            .O(N__23298),
            .I(\QuadInstance2.delayedCh_BZ0Z_0 ));
    InMux I__4183 (
            .O(N__23295),
            .I(N__23292));
    LocalMux I__4182 (
            .O(N__23292),
            .I(N__23289));
    Span4Mux_h I__4181 (
            .O(N__23289),
            .I(N__23286));
    Span4Mux_h I__4180 (
            .O(N__23286),
            .I(N__23283));
    Odrv4 I__4179 (
            .O(N__23283),
            .I(ch4_B_c));
    InMux I__4178 (
            .O(N__23280),
            .I(N__23277));
    LocalMux I__4177 (
            .O(N__23277),
            .I(N__23274));
    Span4Mux_h I__4176 (
            .O(N__23274),
            .I(N__23271));
    Span4Mux_h I__4175 (
            .O(N__23271),
            .I(N__23268));
    Odrv4 I__4174 (
            .O(N__23268),
            .I(ch4_A_c));
    CascadeMux I__4173 (
            .O(N__23265),
            .I(N__23260));
    InMux I__4172 (
            .O(N__23264),
            .I(N__23257));
    InMux I__4171 (
            .O(N__23263),
            .I(N__23254));
    InMux I__4170 (
            .O(N__23260),
            .I(N__23251));
    LocalMux I__4169 (
            .O(N__23257),
            .I(N__23246));
    LocalMux I__4168 (
            .O(N__23254),
            .I(N__23246));
    LocalMux I__4167 (
            .O(N__23251),
            .I(dataRead1_4));
    Odrv4 I__4166 (
            .O(N__23246),
            .I(dataRead1_4));
    CascadeMux I__4165 (
            .O(N__23241),
            .I(N__23238));
    InMux I__4164 (
            .O(N__23238),
            .I(N__23235));
    LocalMux I__4163 (
            .O(N__23235),
            .I(\QuadInstance1.Quad_RNIRK0OZ0Z_4 ));
    InMux I__4162 (
            .O(N__23232),
            .I(N__23228));
    InMux I__4161 (
            .O(N__23231),
            .I(N__23225));
    LocalMux I__4160 (
            .O(N__23228),
            .I(N__23222));
    LocalMux I__4159 (
            .O(N__23225),
            .I(\QuadInstance1.delayedCh_BZ0Z_1 ));
    Odrv4 I__4158 (
            .O(N__23222),
            .I(\QuadInstance1.delayedCh_BZ0Z_1 ));
    CascadeMux I__4157 (
            .O(N__23217),
            .I(\PWMInstance4.un1_periodCounter12_1_0_a2_0_0_cascade_ ));
    InMux I__4156 (
            .O(N__23214),
            .I(N__23211));
    LocalMux I__4155 (
            .O(N__23211),
            .I(\PWMInstance4.PWMPulseWidthCountZ0Z_4 ));
    InMux I__4154 (
            .O(N__23208),
            .I(N__23205));
    LocalMux I__4153 (
            .O(N__23205),
            .I(\PWMInstance4.PWMPulseWidthCountZ0Z_5 ));
    InMux I__4152 (
            .O(N__23202),
            .I(N__23199));
    LocalMux I__4151 (
            .O(N__23199),
            .I(\PWMInstance4.PWMPulseWidthCountZ0Z_10 ));
    InMux I__4150 (
            .O(N__23196),
            .I(N__23192));
    InMux I__4149 (
            .O(N__23195),
            .I(N__23189));
    LocalMux I__4148 (
            .O(N__23192),
            .I(N__23183));
    LocalMux I__4147 (
            .O(N__23189),
            .I(N__23183));
    InMux I__4146 (
            .O(N__23188),
            .I(N__23180));
    Odrv4 I__4145 (
            .O(N__23183),
            .I(\PWMInstance6.periodCounterZ0Z_15 ));
    LocalMux I__4144 (
            .O(N__23180),
            .I(\PWMInstance6.periodCounterZ0Z_15 ));
    InMux I__4143 (
            .O(N__23175),
            .I(N__23171));
    InMux I__4142 (
            .O(N__23174),
            .I(N__23168));
    LocalMux I__4141 (
            .O(N__23171),
            .I(N__23162));
    LocalMux I__4140 (
            .O(N__23168),
            .I(N__23162));
    InMux I__4139 (
            .O(N__23167),
            .I(N__23159));
    Odrv4 I__4138 (
            .O(N__23162),
            .I(\PWMInstance6.periodCounterZ0Z_14 ));
    LocalMux I__4137 (
            .O(N__23159),
            .I(\PWMInstance6.periodCounterZ0Z_14 ));
    CascadeMux I__4136 (
            .O(N__23154),
            .I(N__23151));
    InMux I__4135 (
            .O(N__23151),
            .I(N__23148));
    LocalMux I__4134 (
            .O(N__23148),
            .I(\PWMInstance6.un1_PWMPulseWidthCount_0_I_21_c_RNO_5 ));
    InMux I__4133 (
            .O(N__23145),
            .I(N__23142));
    LocalMux I__4132 (
            .O(N__23142),
            .I(\PWMInstance6.PWMPulseWidthCountZ0Z_14 ));
    CascadeMux I__4131 (
            .O(N__23139),
            .I(N__23136));
    InMux I__4130 (
            .O(N__23136),
            .I(N__23133));
    LocalMux I__4129 (
            .O(N__23133),
            .I(\PWMInstance6.PWMPulseWidthCountZ0Z_15 ));
    InMux I__4128 (
            .O(N__23130),
            .I(N__23125));
    InMux I__4127 (
            .O(N__23129),
            .I(N__23122));
    InMux I__4126 (
            .O(N__23128),
            .I(N__23119));
    LocalMux I__4125 (
            .O(N__23125),
            .I(N__23116));
    LocalMux I__4124 (
            .O(N__23122),
            .I(\PWMInstance6.periodCounterZ0Z_10 ));
    LocalMux I__4123 (
            .O(N__23119),
            .I(\PWMInstance6.periodCounterZ0Z_10 ));
    Odrv12 I__4122 (
            .O(N__23116),
            .I(\PWMInstance6.periodCounterZ0Z_10 ));
    InMux I__4121 (
            .O(N__23109),
            .I(N__23106));
    LocalMux I__4120 (
            .O(N__23106),
            .I(\PWMInstance6.PWMPulseWidthCountZ0Z_11 ));
    CascadeMux I__4119 (
            .O(N__23103),
            .I(N__23099));
    CascadeMux I__4118 (
            .O(N__23102),
            .I(N__23095));
    InMux I__4117 (
            .O(N__23099),
            .I(N__23092));
    InMux I__4116 (
            .O(N__23098),
            .I(N__23089));
    InMux I__4115 (
            .O(N__23095),
            .I(N__23086));
    LocalMux I__4114 (
            .O(N__23092),
            .I(N__23083));
    LocalMux I__4113 (
            .O(N__23089),
            .I(\PWMInstance6.periodCounterZ0Z_11 ));
    LocalMux I__4112 (
            .O(N__23086),
            .I(\PWMInstance6.periodCounterZ0Z_11 ));
    Odrv4 I__4111 (
            .O(N__23083),
            .I(\PWMInstance6.periodCounterZ0Z_11 ));
    CascadeMux I__4110 (
            .O(N__23076),
            .I(N__23073));
    InMux I__4109 (
            .O(N__23073),
            .I(N__23070));
    LocalMux I__4108 (
            .O(N__23070),
            .I(\PWMInstance6.un1_PWMPulseWidthCount_0_I_33_c_RNO_5 ));
    InMux I__4107 (
            .O(N__23067),
            .I(N__23064));
    LocalMux I__4106 (
            .O(N__23064),
            .I(\PWMInstance6.PWMPulseWidthCountZ0Z_10 ));
    InMux I__4105 (
            .O(N__23061),
            .I(N__23058));
    LocalMux I__4104 (
            .O(N__23058),
            .I(\PWMInstance6.PWMPulseWidthCountZ0Z_13 ));
    InMux I__4103 (
            .O(N__23055),
            .I(N__23050));
    InMux I__4102 (
            .O(N__23054),
            .I(N__23047));
    InMux I__4101 (
            .O(N__23053),
            .I(N__23044));
    LocalMux I__4100 (
            .O(N__23050),
            .I(N__23041));
    LocalMux I__4099 (
            .O(N__23047),
            .I(\PWMInstance6.periodCounterZ0Z_12 ));
    LocalMux I__4098 (
            .O(N__23044),
            .I(\PWMInstance6.periodCounterZ0Z_12 ));
    Odrv4 I__4097 (
            .O(N__23041),
            .I(\PWMInstance6.periodCounterZ0Z_12 ));
    CascadeMux I__4096 (
            .O(N__23034),
            .I(N__23031));
    InMux I__4095 (
            .O(N__23031),
            .I(N__23027));
    InMux I__4094 (
            .O(N__23030),
            .I(N__23023));
    LocalMux I__4093 (
            .O(N__23027),
            .I(N__23020));
    InMux I__4092 (
            .O(N__23026),
            .I(N__23017));
    LocalMux I__4091 (
            .O(N__23023),
            .I(\PWMInstance6.periodCounterZ0Z_13 ));
    Odrv4 I__4090 (
            .O(N__23020),
            .I(\PWMInstance6.periodCounterZ0Z_13 ));
    LocalMux I__4089 (
            .O(N__23017),
            .I(\PWMInstance6.periodCounterZ0Z_13 ));
    InMux I__4088 (
            .O(N__23010),
            .I(N__23007));
    LocalMux I__4087 (
            .O(N__23007),
            .I(\PWMInstance6.PWMPulseWidthCountZ0Z_12 ));
    InMux I__4086 (
            .O(N__23004),
            .I(N__23001));
    LocalMux I__4085 (
            .O(N__23001),
            .I(\PWMInstance6.un1_PWMPulseWidthCount_0_I_39_c_RNO_5 ));
    CascadeMux I__4084 (
            .O(N__22998),
            .I(data_received_esr_RNIMIH31Z0Z_19_cascade_));
    InMux I__4083 (
            .O(N__22995),
            .I(N__22990));
    InMux I__4082 (
            .O(N__22994),
            .I(N__22985));
    InMux I__4081 (
            .O(N__22993),
            .I(N__22985));
    LocalMux I__4080 (
            .O(N__22990),
            .I(data_receivedZ0Z_19));
    LocalMux I__4079 (
            .O(N__22985),
            .I(data_receivedZ0Z_19));
    CascadeMux I__4078 (
            .O(N__22980),
            .I(N__22975));
    CascadeMux I__4077 (
            .O(N__22979),
            .I(N__22972));
    InMux I__4076 (
            .O(N__22978),
            .I(N__22965));
    InMux I__4075 (
            .O(N__22975),
            .I(N__22965));
    InMux I__4074 (
            .O(N__22972),
            .I(N__22965));
    LocalMux I__4073 (
            .O(N__22965),
            .I(data_receivedZ0Z_23));
    CascadeMux I__4072 (
            .O(N__22962),
            .I(data_received_esr_RNIMIH31_0Z0Z_19_cascade_));
    InMux I__4071 (
            .O(N__22959),
            .I(N__22956));
    LocalMux I__4070 (
            .O(N__22956),
            .I(N__22953));
    Span4Mux_h I__4069 (
            .O(N__22953),
            .I(N__22950));
    Odrv4 I__4068 (
            .O(N__22950),
            .I(\PWMInstance6.PWMPulseWidthCountZ0Z_5 ));
    InMux I__4067 (
            .O(N__22947),
            .I(N__22944));
    LocalMux I__4066 (
            .O(N__22944),
            .I(\PWMInstance6.PWMPulseWidthCountZ0Z_8 ));
    InMux I__4065 (
            .O(N__22941),
            .I(N__22938));
    LocalMux I__4064 (
            .O(N__22938),
            .I(N__22935));
    Odrv4 I__4063 (
            .O(N__22935),
            .I(OutRegZ0Z_11));
    CascadeMux I__4062 (
            .O(N__22932),
            .I(OutReg_esr_RNO_0Z0Z_12_cascade_));
    InMux I__4061 (
            .O(N__22929),
            .I(N__22926));
    LocalMux I__4060 (
            .O(N__22926),
            .I(OutRegZ0Z_12));
    InMux I__4059 (
            .O(N__22923),
            .I(N__22919));
    InMux I__4058 (
            .O(N__22922),
            .I(N__22916));
    LocalMux I__4057 (
            .O(N__22919),
            .I(data_receivedZ0Z_12));
    LocalMux I__4056 (
            .O(N__22916),
            .I(data_receivedZ0Z_12));
    InMux I__4055 (
            .O(N__22911),
            .I(N__22907));
    InMux I__4054 (
            .O(N__22910),
            .I(N__22904));
    LocalMux I__4053 (
            .O(N__22907),
            .I(data_receivedZ0Z_13));
    LocalMux I__4052 (
            .O(N__22904),
            .I(data_receivedZ0Z_13));
    InMux I__4051 (
            .O(N__22899),
            .I(N__22895));
    InMux I__4050 (
            .O(N__22898),
            .I(N__22892));
    LocalMux I__4049 (
            .O(N__22895),
            .I(data_receivedZ0Z_14));
    LocalMux I__4048 (
            .O(N__22892),
            .I(data_receivedZ0Z_14));
    InMux I__4047 (
            .O(N__22887),
            .I(N__22883));
    InMux I__4046 (
            .O(N__22886),
            .I(N__22880));
    LocalMux I__4045 (
            .O(N__22883),
            .I(data_receivedZ0Z_10));
    LocalMux I__4044 (
            .O(N__22880),
            .I(data_receivedZ0Z_10));
    InMux I__4043 (
            .O(N__22875),
            .I(N__22871));
    InMux I__4042 (
            .O(N__22874),
            .I(N__22868));
    LocalMux I__4041 (
            .O(N__22871),
            .I(data_receivedZ0Z_11));
    LocalMux I__4040 (
            .O(N__22868),
            .I(data_receivedZ0Z_11));
    InMux I__4039 (
            .O(N__22863),
            .I(N__22858));
    InMux I__4038 (
            .O(N__22862),
            .I(N__22855));
    InMux I__4037 (
            .O(N__22861),
            .I(N__22852));
    LocalMux I__4036 (
            .O(N__22858),
            .I(\QuadInstance6.delayedCh_AZ0Z_1 ));
    LocalMux I__4035 (
            .O(N__22855),
            .I(\QuadInstance6.delayedCh_AZ0Z_1 ));
    LocalMux I__4034 (
            .O(N__22852),
            .I(\QuadInstance6.delayedCh_AZ0Z_1 ));
    InMux I__4033 (
            .O(N__22845),
            .I(N__22842));
    LocalMux I__4032 (
            .O(N__22842),
            .I(\QuadInstance6.delayedCh_AZ0Z_2 ));
    CascadeMux I__4031 (
            .O(N__22839),
            .I(N__22835));
    InMux I__4030 (
            .O(N__22838),
            .I(N__22832));
    InMux I__4029 (
            .O(N__22835),
            .I(N__22829));
    LocalMux I__4028 (
            .O(N__22832),
            .I(N__22826));
    LocalMux I__4027 (
            .O(N__22829),
            .I(N__22823));
    Span4Mux_v I__4026 (
            .O(N__22826),
            .I(N__22819));
    Span4Mux_h I__4025 (
            .O(N__22823),
            .I(N__22816));
    InMux I__4024 (
            .O(N__22822),
            .I(N__22813));
    Odrv4 I__4023 (
            .O(N__22819),
            .I(dataRead6_13));
    Odrv4 I__4022 (
            .O(N__22816),
            .I(dataRead6_13));
    LocalMux I__4021 (
            .O(N__22813),
            .I(dataRead6_13));
    InMux I__4020 (
            .O(N__22806),
            .I(N__22802));
    CascadeMux I__4019 (
            .O(N__22805),
            .I(N__22799));
    LocalMux I__4018 (
            .O(N__22802),
            .I(N__22784));
    InMux I__4017 (
            .O(N__22799),
            .I(N__22780));
    InMux I__4016 (
            .O(N__22798),
            .I(N__22777));
    InMux I__4015 (
            .O(N__22797),
            .I(N__22772));
    InMux I__4014 (
            .O(N__22796),
            .I(N__22772));
    InMux I__4013 (
            .O(N__22795),
            .I(N__22765));
    InMux I__4012 (
            .O(N__22794),
            .I(N__22765));
    InMux I__4011 (
            .O(N__22793),
            .I(N__22765));
    InMux I__4010 (
            .O(N__22792),
            .I(N__22762));
    InMux I__4009 (
            .O(N__22791),
            .I(N__22759));
    InMux I__4008 (
            .O(N__22790),
            .I(N__22750));
    InMux I__4007 (
            .O(N__22789),
            .I(N__22743));
    InMux I__4006 (
            .O(N__22788),
            .I(N__22743));
    InMux I__4005 (
            .O(N__22787),
            .I(N__22743));
    Span4Mux_v I__4004 (
            .O(N__22784),
            .I(N__22740));
    InMux I__4003 (
            .O(N__22783),
            .I(N__22737));
    LocalMux I__4002 (
            .O(N__22780),
            .I(N__22730));
    LocalMux I__4001 (
            .O(N__22777),
            .I(N__22730));
    LocalMux I__4000 (
            .O(N__22772),
            .I(N__22730));
    LocalMux I__3999 (
            .O(N__22765),
            .I(N__22723));
    LocalMux I__3998 (
            .O(N__22762),
            .I(N__22723));
    LocalMux I__3997 (
            .O(N__22759),
            .I(N__22723));
    CascadeMux I__3996 (
            .O(N__22758),
            .I(N__22714));
    CascadeMux I__3995 (
            .O(N__22757),
            .I(N__22711));
    CascadeMux I__3994 (
            .O(N__22756),
            .I(N__22707));
    InMux I__3993 (
            .O(N__22755),
            .I(N__22701));
    InMux I__3992 (
            .O(N__22754),
            .I(N__22698));
    InMux I__3991 (
            .O(N__22753),
            .I(N__22695));
    LocalMux I__3990 (
            .O(N__22750),
            .I(N__22688));
    LocalMux I__3989 (
            .O(N__22743),
            .I(N__22688));
    Span4Mux_h I__3988 (
            .O(N__22740),
            .I(N__22688));
    LocalMux I__3987 (
            .O(N__22737),
            .I(N__22681));
    Sp12to4 I__3986 (
            .O(N__22730),
            .I(N__22681));
    Span12Mux_s3_v I__3985 (
            .O(N__22723),
            .I(N__22681));
    InMux I__3984 (
            .O(N__22722),
            .I(N__22676));
    InMux I__3983 (
            .O(N__22721),
            .I(N__22676));
    InMux I__3982 (
            .O(N__22720),
            .I(N__22667));
    InMux I__3981 (
            .O(N__22719),
            .I(N__22667));
    InMux I__3980 (
            .O(N__22718),
            .I(N__22667));
    InMux I__3979 (
            .O(N__22717),
            .I(N__22667));
    InMux I__3978 (
            .O(N__22714),
            .I(N__22652));
    InMux I__3977 (
            .O(N__22711),
            .I(N__22652));
    InMux I__3976 (
            .O(N__22710),
            .I(N__22652));
    InMux I__3975 (
            .O(N__22707),
            .I(N__22652));
    InMux I__3974 (
            .O(N__22706),
            .I(N__22652));
    InMux I__3973 (
            .O(N__22705),
            .I(N__22652));
    InMux I__3972 (
            .O(N__22704),
            .I(N__22652));
    LocalMux I__3971 (
            .O(N__22701),
            .I(quadWriteZ0Z_6));
    LocalMux I__3970 (
            .O(N__22698),
            .I(quadWriteZ0Z_6));
    LocalMux I__3969 (
            .O(N__22695),
            .I(quadWriteZ0Z_6));
    Odrv4 I__3968 (
            .O(N__22688),
            .I(quadWriteZ0Z_6));
    Odrv12 I__3967 (
            .O(N__22681),
            .I(quadWriteZ0Z_6));
    LocalMux I__3966 (
            .O(N__22676),
            .I(quadWriteZ0Z_6));
    LocalMux I__3965 (
            .O(N__22667),
            .I(quadWriteZ0Z_6));
    LocalMux I__3964 (
            .O(N__22652),
            .I(quadWriteZ0Z_6));
    InMux I__3963 (
            .O(N__22635),
            .I(N__22627));
    InMux I__3962 (
            .O(N__22634),
            .I(N__22624));
    CascadeMux I__3961 (
            .O(N__22633),
            .I(N__22621));
    CascadeMux I__3960 (
            .O(N__22632),
            .I(N__22618));
    CascadeMux I__3959 (
            .O(N__22631),
            .I(N__22615));
    CascadeMux I__3958 (
            .O(N__22630),
            .I(N__22611));
    LocalMux I__3957 (
            .O(N__22627),
            .I(N__22599));
    LocalMux I__3956 (
            .O(N__22624),
            .I(N__22599));
    InMux I__3955 (
            .O(N__22621),
            .I(N__22594));
    InMux I__3954 (
            .O(N__22618),
            .I(N__22594));
    InMux I__3953 (
            .O(N__22615),
            .I(N__22587));
    InMux I__3952 (
            .O(N__22614),
            .I(N__22587));
    InMux I__3951 (
            .O(N__22611),
            .I(N__22587));
    InMux I__3950 (
            .O(N__22610),
            .I(N__22572));
    InMux I__3949 (
            .O(N__22609),
            .I(N__22572));
    InMux I__3948 (
            .O(N__22608),
            .I(N__22572));
    InMux I__3947 (
            .O(N__22607),
            .I(N__22572));
    InMux I__3946 (
            .O(N__22606),
            .I(N__22572));
    InMux I__3945 (
            .O(N__22605),
            .I(N__22572));
    InMux I__3944 (
            .O(N__22604),
            .I(N__22572));
    Odrv12 I__3943 (
            .O(N__22599),
            .I(\QuadInstance6.un1_count_enable_i_a2_0_1 ));
    LocalMux I__3942 (
            .O(N__22594),
            .I(\QuadInstance6.un1_count_enable_i_a2_0_1 ));
    LocalMux I__3941 (
            .O(N__22587),
            .I(\QuadInstance6.un1_count_enable_i_a2_0_1 ));
    LocalMux I__3940 (
            .O(N__22572),
            .I(\QuadInstance6.un1_count_enable_i_a2_0_1 ));
    InMux I__3939 (
            .O(N__22563),
            .I(N__22559));
    InMux I__3938 (
            .O(N__22562),
            .I(N__22556));
    LocalMux I__3937 (
            .O(N__22559),
            .I(N__22543));
    LocalMux I__3936 (
            .O(N__22556),
            .I(N__22543));
    InMux I__3935 (
            .O(N__22555),
            .I(N__22540));
    CascadeMux I__3934 (
            .O(N__22554),
            .I(N__22535));
    CascadeMux I__3933 (
            .O(N__22553),
            .I(N__22530));
    CascadeMux I__3932 (
            .O(N__22552),
            .I(N__22525));
    CascadeMux I__3931 (
            .O(N__22551),
            .I(N__22522));
    InMux I__3930 (
            .O(N__22550),
            .I(N__22519));
    InMux I__3929 (
            .O(N__22549),
            .I(N__22514));
    InMux I__3928 (
            .O(N__22548),
            .I(N__22514));
    Span4Mux_s3_v I__3927 (
            .O(N__22543),
            .I(N__22509));
    LocalMux I__3926 (
            .O(N__22540),
            .I(N__22509));
    InMux I__3925 (
            .O(N__22539),
            .I(N__22500));
    InMux I__3924 (
            .O(N__22538),
            .I(N__22500));
    InMux I__3923 (
            .O(N__22535),
            .I(N__22500));
    InMux I__3922 (
            .O(N__22534),
            .I(N__22500));
    InMux I__3921 (
            .O(N__22533),
            .I(N__22487));
    InMux I__3920 (
            .O(N__22530),
            .I(N__22487));
    InMux I__3919 (
            .O(N__22529),
            .I(N__22487));
    InMux I__3918 (
            .O(N__22528),
            .I(N__22487));
    InMux I__3917 (
            .O(N__22525),
            .I(N__22487));
    InMux I__3916 (
            .O(N__22522),
            .I(N__22487));
    LocalMux I__3915 (
            .O(N__22519),
            .I(\QuadInstance6.count_enable ));
    LocalMux I__3914 (
            .O(N__22514),
            .I(\QuadInstance6.count_enable ));
    Odrv4 I__3913 (
            .O(N__22509),
            .I(\QuadInstance6.count_enable ));
    LocalMux I__3912 (
            .O(N__22500),
            .I(\QuadInstance6.count_enable ));
    LocalMux I__3911 (
            .O(N__22487),
            .I(\QuadInstance6.count_enable ));
    InMux I__3910 (
            .O(N__22476),
            .I(N__22473));
    LocalMux I__3909 (
            .O(N__22473),
            .I(N__22470));
    Odrv4 I__3908 (
            .O(N__22470),
            .I(\QuadInstance6.Quad_RNIJHNB1Z0Z_13 ));
    InMux I__3907 (
            .O(N__22467),
            .I(N__22463));
    InMux I__3906 (
            .O(N__22466),
            .I(N__22460));
    LocalMux I__3905 (
            .O(N__22463),
            .I(\QuadInstance6.delayedCh_BZ0Z_1 ));
    LocalMux I__3904 (
            .O(N__22460),
            .I(\QuadInstance6.delayedCh_BZ0Z_1 ));
    InMux I__3903 (
            .O(N__22455),
            .I(N__22452));
    LocalMux I__3902 (
            .O(N__22452),
            .I(N__22447));
    InMux I__3901 (
            .O(N__22451),
            .I(N__22444));
    InMux I__3900 (
            .O(N__22450),
            .I(N__22441));
    Span4Mux_v I__3899 (
            .O(N__22447),
            .I(N__22436));
    LocalMux I__3898 (
            .O(N__22444),
            .I(N__22436));
    LocalMux I__3897 (
            .O(N__22441),
            .I(N__22433));
    Span4Mux_h I__3896 (
            .O(N__22436),
            .I(N__22430));
    Span12Mux_h I__3895 (
            .O(N__22433),
            .I(N__22427));
    Odrv4 I__3894 (
            .O(N__22430),
            .I(dataRead2_11));
    Odrv12 I__3893 (
            .O(N__22427),
            .I(dataRead2_11));
    InMux I__3892 (
            .O(N__22422),
            .I(N__22419));
    LocalMux I__3891 (
            .O(N__22419),
            .I(N__22415));
    InMux I__3890 (
            .O(N__22418),
            .I(N__22411));
    Span4Mux_v I__3889 (
            .O(N__22415),
            .I(N__22408));
    InMux I__3888 (
            .O(N__22414),
            .I(N__22405));
    LocalMux I__3887 (
            .O(N__22411),
            .I(N__22402));
    Odrv4 I__3886 (
            .O(N__22408),
            .I(dataRead3_11));
    LocalMux I__3885 (
            .O(N__22405),
            .I(dataRead3_11));
    Odrv4 I__3884 (
            .O(N__22402),
            .I(dataRead3_11));
    InMux I__3883 (
            .O(N__22395),
            .I(N__22392));
    LocalMux I__3882 (
            .O(N__22392),
            .I(OutReg_0_4_i_m3_i_m3_ns_1_11));
    CascadeMux I__3881 (
            .O(N__22389),
            .I(N__22386));
    InMux I__3880 (
            .O(N__22386),
            .I(N__22382));
    CascadeMux I__3879 (
            .O(N__22385),
            .I(N__22379));
    LocalMux I__3878 (
            .O(N__22382),
            .I(N__22375));
    InMux I__3877 (
            .O(N__22379),
            .I(N__22372));
    InMux I__3876 (
            .O(N__22378),
            .I(N__22369));
    Span4Mux_h I__3875 (
            .O(N__22375),
            .I(N__22366));
    LocalMux I__3874 (
            .O(N__22372),
            .I(dataRead5_12));
    LocalMux I__3873 (
            .O(N__22369),
            .I(dataRead5_12));
    Odrv4 I__3872 (
            .O(N__22366),
            .I(dataRead5_12));
    InMux I__3871 (
            .O(N__22359),
            .I(N__22356));
    LocalMux I__3870 (
            .O(N__22356),
            .I(N__22353));
    Span4Mux_h I__3869 (
            .O(N__22353),
            .I(N__22348));
    InMux I__3868 (
            .O(N__22352),
            .I(N__22345));
    InMux I__3867 (
            .O(N__22351),
            .I(N__22342));
    Span4Mux_h I__3866 (
            .O(N__22348),
            .I(N__22339));
    LocalMux I__3865 (
            .O(N__22345),
            .I(dataRead2_12));
    LocalMux I__3864 (
            .O(N__22342),
            .I(dataRead2_12));
    Odrv4 I__3863 (
            .O(N__22339),
            .I(dataRead2_12));
    CascadeMux I__3862 (
            .O(N__22332),
            .I(N__22328));
    CascadeMux I__3861 (
            .O(N__22331),
            .I(N__22325));
    InMux I__3860 (
            .O(N__22328),
            .I(N__22322));
    InMux I__3859 (
            .O(N__22325),
            .I(N__22319));
    LocalMux I__3858 (
            .O(N__22322),
            .I(N__22316));
    LocalMux I__3857 (
            .O(N__22319),
            .I(N__22312));
    Span4Mux_v I__3856 (
            .O(N__22316),
            .I(N__22309));
    InMux I__3855 (
            .O(N__22315),
            .I(N__22306));
    Span4Mux_h I__3854 (
            .O(N__22312),
            .I(N__22303));
    Span4Mux_h I__3853 (
            .O(N__22309),
            .I(N__22298));
    LocalMux I__3852 (
            .O(N__22306),
            .I(N__22298));
    Odrv4 I__3851 (
            .O(N__22303),
            .I(dataRead3_12));
    Odrv4 I__3850 (
            .O(N__22298),
            .I(dataRead3_12));
    InMux I__3849 (
            .O(N__22293),
            .I(N__22290));
    LocalMux I__3848 (
            .O(N__22290),
            .I(N__22286));
    InMux I__3847 (
            .O(N__22289),
            .I(N__22283));
    Span4Mux_h I__3846 (
            .O(N__22286),
            .I(N__22279));
    LocalMux I__3845 (
            .O(N__22283),
            .I(N__22276));
    InMux I__3844 (
            .O(N__22282),
            .I(N__22273));
    Span4Mux_v I__3843 (
            .O(N__22279),
            .I(N__22268));
    Span4Mux_h I__3842 (
            .O(N__22276),
            .I(N__22268));
    LocalMux I__3841 (
            .O(N__22273),
            .I(dataRead6_12));
    Odrv4 I__3840 (
            .O(N__22268),
            .I(dataRead6_12));
    InMux I__3839 (
            .O(N__22263),
            .I(N__22259));
    InMux I__3838 (
            .O(N__22262),
            .I(N__22256));
    LocalMux I__3837 (
            .O(N__22259),
            .I(N__22253));
    LocalMux I__3836 (
            .O(N__22256),
            .I(N__22249));
    Span4Mux_v I__3835 (
            .O(N__22253),
            .I(N__22246));
    InMux I__3834 (
            .O(N__22252),
            .I(N__22243));
    Span4Mux_v I__3833 (
            .O(N__22249),
            .I(N__22236));
    Span4Mux_h I__3832 (
            .O(N__22246),
            .I(N__22236));
    LocalMux I__3831 (
            .O(N__22243),
            .I(N__22236));
    Odrv4 I__3830 (
            .O(N__22236),
            .I(dataRead7_12));
    CascadeMux I__3829 (
            .O(N__22233),
            .I(OutReg_0_4_i_m3_ns_1_12_cascade_));
    CascadeMux I__3828 (
            .O(N__22230),
            .I(OutReg_esr_RNO_1Z0Z_12_cascade_));
    InMux I__3827 (
            .O(N__22227),
            .I(N__22224));
    LocalMux I__3826 (
            .O(N__22224),
            .I(OutReg_esr_RNO_2Z0Z_12));
    InMux I__3825 (
            .O(N__22221),
            .I(N__22218));
    LocalMux I__3824 (
            .O(N__22218),
            .I(N__22215));
    Span4Mux_v I__3823 (
            .O(N__22215),
            .I(N__22212));
    Odrv4 I__3822 (
            .O(N__22212),
            .I(\QuadInstance6.Quad_RNO_0_6_9 ));
    InMux I__3821 (
            .O(N__22209),
            .I(N__22206));
    LocalMux I__3820 (
            .O(N__22206),
            .I(N__22203));
    Span4Mux_h I__3819 (
            .O(N__22203),
            .I(N__22200));
    Span4Mux_h I__3818 (
            .O(N__22200),
            .I(N__22197));
    Odrv4 I__3817 (
            .O(N__22197),
            .I(\QuadInstance2.Quad_RNO_0_1_1 ));
    InMux I__3816 (
            .O(N__22194),
            .I(N__22178));
    InMux I__3815 (
            .O(N__22193),
            .I(N__22178));
    InMux I__3814 (
            .O(N__22192),
            .I(N__22178));
    InMux I__3813 (
            .O(N__22191),
            .I(N__22175));
    CascadeMux I__3812 (
            .O(N__22190),
            .I(N__22172));
    InMux I__3811 (
            .O(N__22189),
            .I(N__22168));
    InMux I__3810 (
            .O(N__22188),
            .I(N__22165));
    InMux I__3809 (
            .O(N__22187),
            .I(N__22160));
    InMux I__3808 (
            .O(N__22186),
            .I(N__22160));
    InMux I__3807 (
            .O(N__22185),
            .I(N__22156));
    LocalMux I__3806 (
            .O(N__22178),
            .I(N__22151));
    LocalMux I__3805 (
            .O(N__22175),
            .I(N__22151));
    InMux I__3804 (
            .O(N__22172),
            .I(N__22147));
    InMux I__3803 (
            .O(N__22171),
            .I(N__22144));
    LocalMux I__3802 (
            .O(N__22168),
            .I(N__22136));
    LocalMux I__3801 (
            .O(N__22165),
            .I(N__22131));
    LocalMux I__3800 (
            .O(N__22160),
            .I(N__22131));
    InMux I__3799 (
            .O(N__22159),
            .I(N__22128));
    LocalMux I__3798 (
            .O(N__22156),
            .I(N__22123));
    Span4Mux_v I__3797 (
            .O(N__22151),
            .I(N__22123));
    InMux I__3796 (
            .O(N__22150),
            .I(N__22120));
    LocalMux I__3795 (
            .O(N__22147),
            .I(N__22117));
    LocalMux I__3794 (
            .O(N__22144),
            .I(N__22114));
    InMux I__3793 (
            .O(N__22143),
            .I(N__22111));
    InMux I__3792 (
            .O(N__22142),
            .I(N__22089));
    InMux I__3791 (
            .O(N__22141),
            .I(N__22089));
    InMux I__3790 (
            .O(N__22140),
            .I(N__22089));
    InMux I__3789 (
            .O(N__22139),
            .I(N__22089));
    Span4Mux_h I__3788 (
            .O(N__22136),
            .I(N__22084));
    Span4Mux_v I__3787 (
            .O(N__22131),
            .I(N__22084));
    LocalMux I__3786 (
            .O(N__22128),
            .I(N__22077));
    Span4Mux_h I__3785 (
            .O(N__22123),
            .I(N__22077));
    LocalMux I__3784 (
            .O(N__22120),
            .I(N__22077));
    Span4Mux_h I__3783 (
            .O(N__22117),
            .I(N__22070));
    Span4Mux_v I__3782 (
            .O(N__22114),
            .I(N__22070));
    LocalMux I__3781 (
            .O(N__22111),
            .I(N__22070));
    InMux I__3780 (
            .O(N__22110),
            .I(N__22059));
    InMux I__3779 (
            .O(N__22109),
            .I(N__22059));
    InMux I__3778 (
            .O(N__22108),
            .I(N__22059));
    InMux I__3777 (
            .O(N__22107),
            .I(N__22059));
    InMux I__3776 (
            .O(N__22106),
            .I(N__22059));
    InMux I__3775 (
            .O(N__22105),
            .I(N__22042));
    InMux I__3774 (
            .O(N__22104),
            .I(N__22042));
    InMux I__3773 (
            .O(N__22103),
            .I(N__22042));
    InMux I__3772 (
            .O(N__22102),
            .I(N__22042));
    InMux I__3771 (
            .O(N__22101),
            .I(N__22042));
    InMux I__3770 (
            .O(N__22100),
            .I(N__22042));
    InMux I__3769 (
            .O(N__22099),
            .I(N__22042));
    InMux I__3768 (
            .O(N__22098),
            .I(N__22042));
    LocalMux I__3767 (
            .O(N__22089),
            .I(quadWriteZ0Z_2));
    Odrv4 I__3766 (
            .O(N__22084),
            .I(quadWriteZ0Z_2));
    Odrv4 I__3765 (
            .O(N__22077),
            .I(quadWriteZ0Z_2));
    Odrv4 I__3764 (
            .O(N__22070),
            .I(quadWriteZ0Z_2));
    LocalMux I__3763 (
            .O(N__22059),
            .I(quadWriteZ0Z_2));
    LocalMux I__3762 (
            .O(N__22042),
            .I(quadWriteZ0Z_2));
    InMux I__3761 (
            .O(N__22029),
            .I(N__22026));
    LocalMux I__3760 (
            .O(N__22026),
            .I(N__22023));
    Odrv4 I__3759 (
            .O(N__22023),
            .I(\QuadInstance3.Quad_RNO_0_2_1 ));
    InMux I__3758 (
            .O(N__22020),
            .I(N__22009));
    InMux I__3757 (
            .O(N__22019),
            .I(N__22005));
    InMux I__3756 (
            .O(N__22018),
            .I(N__21997));
    InMux I__3755 (
            .O(N__22017),
            .I(N__21994));
    InMux I__3754 (
            .O(N__22016),
            .I(N__21991));
    InMux I__3753 (
            .O(N__22015),
            .I(N__21986));
    InMux I__3752 (
            .O(N__22014),
            .I(N__21986));
    InMux I__3751 (
            .O(N__22013),
            .I(N__21980));
    InMux I__3750 (
            .O(N__22012),
            .I(N__21980));
    LocalMux I__3749 (
            .O(N__22009),
            .I(N__21977));
    InMux I__3748 (
            .O(N__22008),
            .I(N__21974));
    LocalMux I__3747 (
            .O(N__22005),
            .I(N__21971));
    InMux I__3746 (
            .O(N__22004),
            .I(N__21958));
    InMux I__3745 (
            .O(N__22003),
            .I(N__21958));
    InMux I__3744 (
            .O(N__22002),
            .I(N__21958));
    InMux I__3743 (
            .O(N__22001),
            .I(N__21958));
    InMux I__3742 (
            .O(N__22000),
            .I(N__21958));
    LocalMux I__3741 (
            .O(N__21997),
            .I(N__21949));
    LocalMux I__3740 (
            .O(N__21994),
            .I(N__21949));
    LocalMux I__3739 (
            .O(N__21991),
            .I(N__21949));
    LocalMux I__3738 (
            .O(N__21986),
            .I(N__21949));
    InMux I__3737 (
            .O(N__21985),
            .I(N__21946));
    LocalMux I__3736 (
            .O(N__21980),
            .I(N__21941));
    Span4Mux_v I__3735 (
            .O(N__21977),
            .I(N__21941));
    LocalMux I__3734 (
            .O(N__21974),
            .I(N__21936));
    Span4Mux_h I__3733 (
            .O(N__21971),
            .I(N__21936));
    CascadeMux I__3732 (
            .O(N__21970),
            .I(N__21930));
    CascadeMux I__3731 (
            .O(N__21969),
            .I(N__21924));
    LocalMux I__3730 (
            .O(N__21958),
            .I(N__21912));
    Span4Mux_v I__3729 (
            .O(N__21949),
            .I(N__21912));
    LocalMux I__3728 (
            .O(N__21946),
            .I(N__21905));
    Span4Mux_h I__3727 (
            .O(N__21941),
            .I(N__21905));
    Span4Mux_v I__3726 (
            .O(N__21936),
            .I(N__21905));
    InMux I__3725 (
            .O(N__21935),
            .I(N__21900));
    InMux I__3724 (
            .O(N__21934),
            .I(N__21900));
    InMux I__3723 (
            .O(N__21933),
            .I(N__21897));
    InMux I__3722 (
            .O(N__21930),
            .I(N__21894));
    InMux I__3721 (
            .O(N__21929),
            .I(N__21881));
    InMux I__3720 (
            .O(N__21928),
            .I(N__21881));
    InMux I__3719 (
            .O(N__21927),
            .I(N__21881));
    InMux I__3718 (
            .O(N__21924),
            .I(N__21881));
    InMux I__3717 (
            .O(N__21923),
            .I(N__21881));
    InMux I__3716 (
            .O(N__21922),
            .I(N__21881));
    InMux I__3715 (
            .O(N__21921),
            .I(N__21870));
    InMux I__3714 (
            .O(N__21920),
            .I(N__21870));
    InMux I__3713 (
            .O(N__21919),
            .I(N__21870));
    InMux I__3712 (
            .O(N__21918),
            .I(N__21870));
    InMux I__3711 (
            .O(N__21917),
            .I(N__21870));
    Odrv4 I__3710 (
            .O(N__21912),
            .I(quadWriteZ0Z_3));
    Odrv4 I__3709 (
            .O(N__21905),
            .I(quadWriteZ0Z_3));
    LocalMux I__3708 (
            .O(N__21900),
            .I(quadWriteZ0Z_3));
    LocalMux I__3707 (
            .O(N__21897),
            .I(quadWriteZ0Z_3));
    LocalMux I__3706 (
            .O(N__21894),
            .I(quadWriteZ0Z_3));
    LocalMux I__3705 (
            .O(N__21881),
            .I(quadWriteZ0Z_3));
    LocalMux I__3704 (
            .O(N__21870),
            .I(quadWriteZ0Z_3));
    InMux I__3703 (
            .O(N__21855),
            .I(N__21852));
    LocalMux I__3702 (
            .O(N__21852),
            .I(N__21849));
    Odrv4 I__3701 (
            .O(N__21849),
            .I(\QuadInstance3.Quad_RNO_0_3_4 ));
    InMux I__3700 (
            .O(N__21846),
            .I(N__21842));
    CascadeMux I__3699 (
            .O(N__21845),
            .I(N__21839));
    LocalMux I__3698 (
            .O(N__21842),
            .I(N__21835));
    InMux I__3697 (
            .O(N__21839),
            .I(N__21832));
    InMux I__3696 (
            .O(N__21838),
            .I(N__21829));
    Span4Mux_h I__3695 (
            .O(N__21835),
            .I(N__21826));
    LocalMux I__3694 (
            .O(N__21832),
            .I(N__21823));
    LocalMux I__3693 (
            .O(N__21829),
            .I(N__21820));
    Odrv4 I__3692 (
            .O(N__21826),
            .I(dataRead3_4));
    Odrv4 I__3691 (
            .O(N__21823),
            .I(dataRead3_4));
    Odrv12 I__3690 (
            .O(N__21820),
            .I(dataRead3_4));
    InMux I__3689 (
            .O(N__21813),
            .I(N__21810));
    LocalMux I__3688 (
            .O(N__21810),
            .I(\QuadInstance1.Quad_RNO_0_1_9 ));
    InMux I__3687 (
            .O(N__21807),
            .I(N__21804));
    LocalMux I__3686 (
            .O(N__21804),
            .I(N__21796));
    CascadeMux I__3685 (
            .O(N__21803),
            .I(N__21788));
    CascadeMux I__3684 (
            .O(N__21802),
            .I(N__21783));
    CascadeMux I__3683 (
            .O(N__21801),
            .I(N__21778));
    CascadeMux I__3682 (
            .O(N__21800),
            .I(N__21774));
    CascadeMux I__3681 (
            .O(N__21799),
            .I(N__21771));
    Span12Mux_s8_v I__3680 (
            .O(N__21796),
            .I(N__21768));
    InMux I__3679 (
            .O(N__21795),
            .I(N__21765));
    InMux I__3678 (
            .O(N__21794),
            .I(N__21758));
    InMux I__3677 (
            .O(N__21793),
            .I(N__21758));
    InMux I__3676 (
            .O(N__21792),
            .I(N__21758));
    InMux I__3675 (
            .O(N__21791),
            .I(N__21755));
    InMux I__3674 (
            .O(N__21788),
            .I(N__21744));
    InMux I__3673 (
            .O(N__21787),
            .I(N__21744));
    InMux I__3672 (
            .O(N__21786),
            .I(N__21744));
    InMux I__3671 (
            .O(N__21783),
            .I(N__21744));
    InMux I__3670 (
            .O(N__21782),
            .I(N__21744));
    InMux I__3669 (
            .O(N__21781),
            .I(N__21733));
    InMux I__3668 (
            .O(N__21778),
            .I(N__21733));
    InMux I__3667 (
            .O(N__21777),
            .I(N__21733));
    InMux I__3666 (
            .O(N__21774),
            .I(N__21733));
    InMux I__3665 (
            .O(N__21771),
            .I(N__21733));
    Odrv12 I__3664 (
            .O(N__21768),
            .I(\QuadInstance7.count_enable ));
    LocalMux I__3663 (
            .O(N__21765),
            .I(\QuadInstance7.count_enable ));
    LocalMux I__3662 (
            .O(N__21758),
            .I(\QuadInstance7.count_enable ));
    LocalMux I__3661 (
            .O(N__21755),
            .I(\QuadInstance7.count_enable ));
    LocalMux I__3660 (
            .O(N__21744),
            .I(\QuadInstance7.count_enable ));
    LocalMux I__3659 (
            .O(N__21733),
            .I(\QuadInstance7.count_enable ));
    CascadeMux I__3658 (
            .O(N__21720),
            .I(N__21716));
    CascadeMux I__3657 (
            .O(N__21719),
            .I(N__21713));
    InMux I__3656 (
            .O(N__21716),
            .I(N__21710));
    InMux I__3655 (
            .O(N__21713),
            .I(N__21707));
    LocalMux I__3654 (
            .O(N__21710),
            .I(\QuadInstance6.delayedCh_BZ0Z_2 ));
    LocalMux I__3653 (
            .O(N__21707),
            .I(\QuadInstance6.delayedCh_BZ0Z_2 ));
    CascadeMux I__3652 (
            .O(N__21702),
            .I(N__21699));
    InMux I__3651 (
            .O(N__21699),
            .I(N__21696));
    LocalMux I__3650 (
            .O(N__21696),
            .I(N__21693));
    Odrv4 I__3649 (
            .O(N__21693),
            .I(\QuadInstance6.Quad_RNIGENB1Z0Z_10 ));
    InMux I__3648 (
            .O(N__21690),
            .I(bfn_13_7_0_));
    InMux I__3647 (
            .O(N__21687),
            .I(\QuadInstance1.un1_Quad_cry_8 ));
    InMux I__3646 (
            .O(N__21684),
            .I(N__21681));
    LocalMux I__3645 (
            .O(N__21681),
            .I(\QuadInstance1.Quad_RNO_0_1_10 ));
    InMux I__3644 (
            .O(N__21678),
            .I(\QuadInstance1.un1_Quad_cry_9 ));
    InMux I__3643 (
            .O(N__21675),
            .I(N__21672));
    LocalMux I__3642 (
            .O(N__21672),
            .I(N__21669));
    Odrv4 I__3641 (
            .O(N__21669),
            .I(\QuadInstance1.Quad_RNO_0_1_11 ));
    InMux I__3640 (
            .O(N__21666),
            .I(\QuadInstance1.un1_Quad_cry_10 ));
    InMux I__3639 (
            .O(N__21663),
            .I(\QuadInstance1.un1_Quad_cry_11 ));
    InMux I__3638 (
            .O(N__21660),
            .I(\QuadInstance1.un1_Quad_cry_12 ));
    InMux I__3637 (
            .O(N__21657),
            .I(N__21654));
    LocalMux I__3636 (
            .O(N__21654),
            .I(\QuadInstance1.Quad_RNO_0_1_14 ));
    InMux I__3635 (
            .O(N__21651),
            .I(\QuadInstance1.un1_Quad_cry_13 ));
    InMux I__3634 (
            .O(N__21648),
            .I(\QuadInstance1.un1_Quad_cry_14 ));
    InMux I__3633 (
            .O(N__21645),
            .I(N__21642));
    LocalMux I__3632 (
            .O(N__21642),
            .I(N__21639));
    Odrv4 I__3631 (
            .O(N__21639),
            .I(\QuadInstance1.Quad_RNO_0_0_1 ));
    InMux I__3630 (
            .O(N__21636),
            .I(\QuadInstance1.un1_Quad_cry_0 ));
    InMux I__3629 (
            .O(N__21633),
            .I(N__21630));
    LocalMux I__3628 (
            .O(N__21630),
            .I(N__21627));
    Span4Mux_h I__3627 (
            .O(N__21627),
            .I(N__21624));
    Span4Mux_h I__3626 (
            .O(N__21624),
            .I(N__21621));
    Odrv4 I__3625 (
            .O(N__21621),
            .I(\QuadInstance1.Quad_RNO_0_1_2 ));
    InMux I__3624 (
            .O(N__21618),
            .I(\QuadInstance1.un1_Quad_cry_1 ));
    InMux I__3623 (
            .O(N__21615),
            .I(N__21612));
    LocalMux I__3622 (
            .O(N__21612),
            .I(N__21609));
    Span4Mux_v I__3621 (
            .O(N__21609),
            .I(N__21606));
    Odrv4 I__3620 (
            .O(N__21606),
            .I(\QuadInstance1.Quad_RNO_0_1_3 ));
    InMux I__3619 (
            .O(N__21603),
            .I(\QuadInstance1.un1_Quad_cry_2 ));
    InMux I__3618 (
            .O(N__21600),
            .I(N__21597));
    LocalMux I__3617 (
            .O(N__21597),
            .I(\QuadInstance1.Quad_RNO_0_1_4 ));
    InMux I__3616 (
            .O(N__21594),
            .I(\QuadInstance1.un1_Quad_cry_3 ));
    InMux I__3615 (
            .O(N__21591),
            .I(N__21588));
    LocalMux I__3614 (
            .O(N__21588),
            .I(N__21585));
    Odrv4 I__3613 (
            .O(N__21585),
            .I(\QuadInstance1.Quad_RNO_0_1_5 ));
    InMux I__3612 (
            .O(N__21582),
            .I(\QuadInstance1.un1_Quad_cry_4 ));
    CascadeMux I__3611 (
            .O(N__21579),
            .I(N__21576));
    InMux I__3610 (
            .O(N__21576),
            .I(N__21573));
    LocalMux I__3609 (
            .O(N__21573),
            .I(N__21570));
    Odrv4 I__3608 (
            .O(N__21570),
            .I(\QuadInstance1.Quad_RNO_0_1_6 ));
    InMux I__3607 (
            .O(N__21567),
            .I(\QuadInstance1.un1_Quad_cry_5 ));
    InMux I__3606 (
            .O(N__21564),
            .I(N__21561));
    LocalMux I__3605 (
            .O(N__21561),
            .I(N__21558));
    Odrv4 I__3604 (
            .O(N__21558),
            .I(\QuadInstance1.Quad_RNO_0_1_7 ));
    InMux I__3603 (
            .O(N__21555),
            .I(\QuadInstance1.un1_Quad_cry_6 ));
    InMux I__3602 (
            .O(N__21552),
            .I(N__21549));
    LocalMux I__3601 (
            .O(N__21549),
            .I(N__21546));
    Span4Mux_v I__3600 (
            .O(N__21546),
            .I(N__21543));
    Odrv4 I__3599 (
            .O(N__21543),
            .I(\QuadInstance1.Quad_RNO_0_1_8 ));
    InMux I__3598 (
            .O(N__21540),
            .I(N__21537));
    LocalMux I__3597 (
            .O(N__21537),
            .I(N__21534));
    Span4Mux_v I__3596 (
            .O(N__21534),
            .I(N__21531));
    Span4Mux_h I__3595 (
            .O(N__21531),
            .I(N__21528));
    Odrv4 I__3594 (
            .O(N__21528),
            .I(ch0_A_c));
    InMux I__3593 (
            .O(N__21525),
            .I(N__21522));
    LocalMux I__3592 (
            .O(N__21522),
            .I(N__21519));
    Span4Mux_h I__3591 (
            .O(N__21519),
            .I(N__21516));
    Odrv4 I__3590 (
            .O(N__21516),
            .I(\QuadInstance3.Quad_RNO_0_3_6 ));
    CascadeMux I__3589 (
            .O(N__21513),
            .I(N__21510));
    InMux I__3588 (
            .O(N__21510),
            .I(N__21507));
    LocalMux I__3587 (
            .O(N__21507),
            .I(\QuadInstance6.Quad_RNO_0_6_4 ));
    InMux I__3586 (
            .O(N__21504),
            .I(N__21501));
    LocalMux I__3585 (
            .O(N__21501),
            .I(N__21497));
    InMux I__3584 (
            .O(N__21500),
            .I(N__21493));
    Span12Mux_v I__3583 (
            .O(N__21497),
            .I(N__21490));
    InMux I__3582 (
            .O(N__21496),
            .I(N__21487));
    LocalMux I__3581 (
            .O(N__21493),
            .I(N__21484));
    Odrv12 I__3580 (
            .O(N__21490),
            .I(dataRead6_4));
    LocalMux I__3579 (
            .O(N__21487),
            .I(dataRead6_4));
    Odrv4 I__3578 (
            .O(N__21484),
            .I(dataRead6_4));
    InMux I__3577 (
            .O(N__21477),
            .I(N__21474));
    LocalMux I__3576 (
            .O(N__21474),
            .I(N__21471));
    Span4Mux_v I__3575 (
            .O(N__21471),
            .I(N__21468));
    Odrv4 I__3574 (
            .O(N__21468),
            .I(\QuadInstance7.Quad_RNO_0_7_4 ));
    InMux I__3573 (
            .O(N__21465),
            .I(N__21461));
    InMux I__3572 (
            .O(N__21464),
            .I(N__21458));
    LocalMux I__3571 (
            .O(N__21461),
            .I(N__21455));
    LocalMux I__3570 (
            .O(N__21458),
            .I(N__21452));
    Span4Mux_v I__3569 (
            .O(N__21455),
            .I(N__21446));
    Span4Mux_v I__3568 (
            .O(N__21452),
            .I(N__21446));
    InMux I__3567 (
            .O(N__21451),
            .I(N__21443));
    Span4Mux_h I__3566 (
            .O(N__21446),
            .I(N__21440));
    LocalMux I__3565 (
            .O(N__21443),
            .I(dataRead7_4));
    Odrv4 I__3564 (
            .O(N__21440),
            .I(dataRead7_4));
    InMux I__3563 (
            .O(N__21435),
            .I(N__21432));
    LocalMux I__3562 (
            .O(N__21432),
            .I(N__21429));
    Odrv12 I__3561 (
            .O(N__21429),
            .I(\PWMInstance6.un1_periodCounter12_1_0_a2_0 ));
    CascadeMux I__3560 (
            .O(N__21426),
            .I(N__21423));
    InMux I__3559 (
            .O(N__21423),
            .I(N__21417));
    InMux I__3558 (
            .O(N__21422),
            .I(N__21414));
    InMux I__3557 (
            .O(N__21421),
            .I(N__21407));
    InMux I__3556 (
            .O(N__21420),
            .I(N__21407));
    LocalMux I__3555 (
            .O(N__21417),
            .I(N__21404));
    LocalMux I__3554 (
            .O(N__21414),
            .I(N__21401));
    InMux I__3553 (
            .O(N__21413),
            .I(N__21398));
    InMux I__3552 (
            .O(N__21412),
            .I(N__21395));
    LocalMux I__3551 (
            .O(N__21407),
            .I(N__21390));
    Span4Mux_v I__3550 (
            .O(N__21404),
            .I(N__21390));
    Odrv4 I__3549 (
            .O(N__21401),
            .I(\PWMInstance6.out_0_sqmuxa ));
    LocalMux I__3548 (
            .O(N__21398),
            .I(\PWMInstance6.out_0_sqmuxa ));
    LocalMux I__3547 (
            .O(N__21395),
            .I(\PWMInstance6.out_0_sqmuxa ));
    Odrv4 I__3546 (
            .O(N__21390),
            .I(\PWMInstance6.out_0_sqmuxa ));
    InMux I__3545 (
            .O(N__21381),
            .I(bfn_12_17_0_));
    IoInMux I__3544 (
            .O(N__21378),
            .I(N__21375));
    LocalMux I__3543 (
            .O(N__21375),
            .I(N__21372));
    Span4Mux_s1_v I__3542 (
            .O(N__21372),
            .I(N__21369));
    Span4Mux_h I__3541 (
            .O(N__21369),
            .I(N__21365));
    InMux I__3540 (
            .O(N__21368),
            .I(N__21362));
    Odrv4 I__3539 (
            .O(N__21365),
            .I(PWM6_c));
    LocalMux I__3538 (
            .O(N__21362),
            .I(PWM6_c));
    IoInMux I__3537 (
            .O(N__21357),
            .I(N__21354));
    LocalMux I__3536 (
            .O(N__21354),
            .I(PWM5_obufLegalizeSB_DFFNet));
    InMux I__3535 (
            .O(N__21351),
            .I(N__21348));
    LocalMux I__3534 (
            .O(N__21348),
            .I(N__21345));
    Span4Mux_h I__3533 (
            .O(N__21345),
            .I(N__21342));
    Odrv4 I__3532 (
            .O(N__21342),
            .I(ch2_A_c));
    InMux I__3531 (
            .O(N__21339),
            .I(N__21336));
    LocalMux I__3530 (
            .O(N__21336),
            .I(N__21333));
    Span12Mux_h I__3529 (
            .O(N__21333),
            .I(N__21330));
    Odrv12 I__3528 (
            .O(N__21330),
            .I(\QuadInstance2.delayedCh_AZ0Z_0 ));
    InMux I__3527 (
            .O(N__21327),
            .I(N__21323));
    InMux I__3526 (
            .O(N__21326),
            .I(N__21320));
    LocalMux I__3525 (
            .O(N__21323),
            .I(N__21317));
    LocalMux I__3524 (
            .O(N__21320),
            .I(N__21313));
    Span4Mux_v I__3523 (
            .O(N__21317),
            .I(N__21310));
    InMux I__3522 (
            .O(N__21316),
            .I(N__21307));
    Odrv12 I__3521 (
            .O(N__21313),
            .I(dataRead5_4));
    Odrv4 I__3520 (
            .O(N__21310),
            .I(dataRead5_4));
    LocalMux I__3519 (
            .O(N__21307),
            .I(dataRead5_4));
    CascadeMux I__3518 (
            .O(N__21300),
            .I(OutReg_ess_RNO_2Z0Z_4_cascade_));
    InMux I__3517 (
            .O(N__21297),
            .I(N__21292));
    InMux I__3516 (
            .O(N__21296),
            .I(N__21289));
    InMux I__3515 (
            .O(N__21295),
            .I(N__21286));
    LocalMux I__3514 (
            .O(N__21292),
            .I(N__21283));
    LocalMux I__3513 (
            .O(N__21289),
            .I(N__21280));
    LocalMux I__3512 (
            .O(N__21286),
            .I(N__21277));
    Span12Mux_s9_h I__3511 (
            .O(N__21283),
            .I(N__21274));
    Span4Mux_h I__3510 (
            .O(N__21280),
            .I(N__21271));
    Span4Mux_v I__3509 (
            .O(N__21277),
            .I(N__21268));
    Odrv12 I__3508 (
            .O(N__21274),
            .I(dataRead2_4));
    Odrv4 I__3507 (
            .O(N__21271),
            .I(dataRead2_4));
    Odrv4 I__3506 (
            .O(N__21268),
            .I(dataRead2_4));
    CascadeMux I__3505 (
            .O(N__21261),
            .I(OutReg_0_4_i_m3_ns_1_4_cascade_));
    InMux I__3504 (
            .O(N__21258),
            .I(N__21255));
    LocalMux I__3503 (
            .O(N__21255),
            .I(OutReg_ess_RNO_1Z0Z_4));
    InMux I__3502 (
            .O(N__21252),
            .I(N__21249));
    LocalMux I__3501 (
            .O(N__21249),
            .I(OutReg_0_5_i_m3_ns_1_4));
    InMux I__3500 (
            .O(N__21246),
            .I(N__21241));
    InMux I__3499 (
            .O(N__21245),
            .I(N__21238));
    InMux I__3498 (
            .O(N__21244),
            .I(N__21235));
    LocalMux I__3497 (
            .O(N__21241),
            .I(\PWMInstance6.periodCounterZ0Z_8 ));
    LocalMux I__3496 (
            .O(N__21238),
            .I(\PWMInstance6.periodCounterZ0Z_8 ));
    LocalMux I__3495 (
            .O(N__21235),
            .I(\PWMInstance6.periodCounterZ0Z_8 ));
    CascadeMux I__3494 (
            .O(N__21228),
            .I(N__21223));
    InMux I__3493 (
            .O(N__21227),
            .I(N__21220));
    InMux I__3492 (
            .O(N__21226),
            .I(N__21217));
    InMux I__3491 (
            .O(N__21223),
            .I(N__21214));
    LocalMux I__3490 (
            .O(N__21220),
            .I(\PWMInstance6.periodCounterZ0Z_9 ));
    LocalMux I__3489 (
            .O(N__21217),
            .I(\PWMInstance6.periodCounterZ0Z_9 ));
    LocalMux I__3488 (
            .O(N__21214),
            .I(\PWMInstance6.periodCounterZ0Z_9 ));
    InMux I__3487 (
            .O(N__21207),
            .I(N__21204));
    LocalMux I__3486 (
            .O(N__21204),
            .I(\PWMInstance6.un1_PWMPulseWidthCount_0_I_1_c_RNO_5 ));
    CascadeMux I__3485 (
            .O(N__21201),
            .I(N__21198));
    InMux I__3484 (
            .O(N__21198),
            .I(N__21195));
    LocalMux I__3483 (
            .O(N__21195),
            .I(N__21192));
    Odrv4 I__3482 (
            .O(N__21192),
            .I(\PWMInstance6.un1_PWMPulseWidthCount_0_I_9_c_RNO_5 ));
    InMux I__3481 (
            .O(N__21189),
            .I(N__21186));
    LocalMux I__3480 (
            .O(N__21186),
            .I(N__21183));
    Odrv4 I__3479 (
            .O(N__21183),
            .I(\PWMInstance6.un1_PWMPulseWidthCount_0_I_15_c_RNO_5 ));
    CascadeMux I__3478 (
            .O(N__21180),
            .I(N__21177));
    InMux I__3477 (
            .O(N__21177),
            .I(N__21174));
    LocalMux I__3476 (
            .O(N__21174),
            .I(\PWMInstance6.un1_PWMPulseWidthCount_0_I_27_c_RNO_5 ));
    InMux I__3475 (
            .O(N__21171),
            .I(N__21168));
    LocalMux I__3474 (
            .O(N__21168),
            .I(\PWMInstance6.un1_PWMPulseWidthCount_0_I_45_c_RNO_5 ));
    CascadeMux I__3473 (
            .O(N__21165),
            .I(\PWMInstance6.un1_periodCounter12_1_0_a2_0_6_cascade_ ));
    CascadeMux I__3472 (
            .O(N__21162),
            .I(N__21159));
    InMux I__3471 (
            .O(N__21159),
            .I(N__21155));
    InMux I__3470 (
            .O(N__21158),
            .I(N__21151));
    LocalMux I__3469 (
            .O(N__21155),
            .I(N__21148));
    InMux I__3468 (
            .O(N__21154),
            .I(N__21145));
    LocalMux I__3467 (
            .O(N__21151),
            .I(\PWMInstance6.periodCounter12 ));
    Odrv4 I__3466 (
            .O(N__21148),
            .I(\PWMInstance6.periodCounter12 ));
    LocalMux I__3465 (
            .O(N__21145),
            .I(\PWMInstance6.periodCounter12 ));
    InMux I__3464 (
            .O(N__21138),
            .I(N__21135));
    LocalMux I__3463 (
            .O(N__21135),
            .I(N__21132));
    Span4Mux_h I__3462 (
            .O(N__21132),
            .I(N__21129));
    Odrv4 I__3461 (
            .O(N__21129),
            .I(\PWMInstance6.un1_periodCounter12_1_0_a2_0_14 ));
    InMux I__3460 (
            .O(N__21126),
            .I(N__21123));
    LocalMux I__3459 (
            .O(N__21123),
            .I(N__21120));
    Span4Mux_v I__3458 (
            .O(N__21120),
            .I(N__21117));
    IoSpan4Mux I__3457 (
            .O(N__21117),
            .I(N__21114));
    Odrv4 I__3456 (
            .O(N__21114),
            .I(ch6_A_c));
    InMux I__3455 (
            .O(N__21111),
            .I(N__21108));
    LocalMux I__3454 (
            .O(N__21108),
            .I(N__21105));
    Span4Mux_v I__3453 (
            .O(N__21105),
            .I(N__21102));
    Odrv4 I__3452 (
            .O(N__21102),
            .I(\QuadInstance6.delayedCh_AZ0Z_0 ));
    InMux I__3451 (
            .O(N__21099),
            .I(N__21096));
    LocalMux I__3450 (
            .O(N__21096),
            .I(N__21093));
    Odrv4 I__3449 (
            .O(N__21093),
            .I(\PWMInstance6.un1_periodCounter12_1_0_a2_0_9 ));
    InMux I__3448 (
            .O(N__21090),
            .I(N__21085));
    InMux I__3447 (
            .O(N__21089),
            .I(N__21080));
    InMux I__3446 (
            .O(N__21088),
            .I(N__21080));
    LocalMux I__3445 (
            .O(N__21085),
            .I(\PWMInstance6.periodCounterZ0Z_0 ));
    LocalMux I__3444 (
            .O(N__21080),
            .I(\PWMInstance6.periodCounterZ0Z_0 ));
    CascadeMux I__3443 (
            .O(N__21075),
            .I(N__21070));
    InMux I__3442 (
            .O(N__21074),
            .I(N__21067));
    InMux I__3441 (
            .O(N__21073),
            .I(N__21064));
    InMux I__3440 (
            .O(N__21070),
            .I(N__21061));
    LocalMux I__3439 (
            .O(N__21067),
            .I(\PWMInstance6.periodCounterZ0Z_1 ));
    LocalMux I__3438 (
            .O(N__21064),
            .I(\PWMInstance6.periodCounterZ0Z_1 ));
    LocalMux I__3437 (
            .O(N__21061),
            .I(\PWMInstance6.periodCounterZ0Z_1 ));
    InMux I__3436 (
            .O(N__21054),
            .I(N__21051));
    LocalMux I__3435 (
            .O(N__21051),
            .I(\PWMInstance6.PWMPulseWidthCountZ0Z_0 ));
    InMux I__3434 (
            .O(N__21048),
            .I(N__21045));
    LocalMux I__3433 (
            .O(N__21045),
            .I(\PWMInstance6.PWMPulseWidthCountZ0Z_1 ));
    CascadeMux I__3432 (
            .O(N__21042),
            .I(N__21038));
    InMux I__3431 (
            .O(N__21041),
            .I(N__21034));
    InMux I__3430 (
            .O(N__21038),
            .I(N__21029));
    InMux I__3429 (
            .O(N__21037),
            .I(N__21029));
    LocalMux I__3428 (
            .O(N__21034),
            .I(\PWMInstance6.periodCounterZ0Z_6 ));
    LocalMux I__3427 (
            .O(N__21029),
            .I(\PWMInstance6.periodCounterZ0Z_6 ));
    InMux I__3426 (
            .O(N__21024),
            .I(N__21019));
    InMux I__3425 (
            .O(N__21023),
            .I(N__21016));
    InMux I__3424 (
            .O(N__21022),
            .I(N__21013));
    LocalMux I__3423 (
            .O(N__21019),
            .I(\PWMInstance6.periodCounterZ0Z_7 ));
    LocalMux I__3422 (
            .O(N__21016),
            .I(\PWMInstance6.periodCounterZ0Z_7 ));
    LocalMux I__3421 (
            .O(N__21013),
            .I(\PWMInstance6.periodCounterZ0Z_7 ));
    InMux I__3420 (
            .O(N__21006),
            .I(N__21003));
    LocalMux I__3419 (
            .O(N__21003),
            .I(\PWMInstance6.PWMPulseWidthCountZ0Z_6 ));
    CascadeMux I__3418 (
            .O(N__21000),
            .I(N__20997));
    InMux I__3417 (
            .O(N__20997),
            .I(N__20994));
    LocalMux I__3416 (
            .O(N__20994),
            .I(\PWMInstance6.PWMPulseWidthCountZ0Z_7 ));
    InMux I__3415 (
            .O(N__20991),
            .I(N__20983));
    InMux I__3414 (
            .O(N__20990),
            .I(N__20983));
    InMux I__3413 (
            .O(N__20989),
            .I(N__20978));
    InMux I__3412 (
            .O(N__20988),
            .I(N__20978));
    LocalMux I__3411 (
            .O(N__20983),
            .I(\PWMInstance6.clkCountZ0Z_0 ));
    LocalMux I__3410 (
            .O(N__20978),
            .I(\PWMInstance6.clkCountZ0Z_0 ));
    CascadeMux I__3409 (
            .O(N__20973),
            .I(N__20970));
    InMux I__3408 (
            .O(N__20970),
            .I(N__20962));
    InMux I__3407 (
            .O(N__20969),
            .I(N__20962));
    InMux I__3406 (
            .O(N__20968),
            .I(N__20957));
    InMux I__3405 (
            .O(N__20967),
            .I(N__20957));
    LocalMux I__3404 (
            .O(N__20962),
            .I(\PWMInstance6.clkCountZ0Z_1 ));
    LocalMux I__3403 (
            .O(N__20957),
            .I(\PWMInstance6.clkCountZ0Z_1 ));
    InMux I__3402 (
            .O(N__20952),
            .I(N__20946));
    InMux I__3401 (
            .O(N__20951),
            .I(N__20946));
    LocalMux I__3400 (
            .O(N__20946),
            .I(pwmWrite_fastZ0Z_6));
    InMux I__3399 (
            .O(N__20943),
            .I(N__20936));
    InMux I__3398 (
            .O(N__20942),
            .I(N__20936));
    InMux I__3397 (
            .O(N__20941),
            .I(N__20933));
    LocalMux I__3396 (
            .O(N__20936),
            .I(pwmWriteZ0Z_6));
    LocalMux I__3395 (
            .O(N__20933),
            .I(pwmWriteZ0Z_6));
    CascadeMux I__3394 (
            .O(N__20928),
            .I(N__20925));
    InMux I__3393 (
            .O(N__20925),
            .I(N__20918));
    InMux I__3392 (
            .O(N__20924),
            .I(N__20918));
    InMux I__3391 (
            .O(N__20923),
            .I(N__20915));
    LocalMux I__3390 (
            .O(N__20918),
            .I(N__20912));
    LocalMux I__3389 (
            .O(N__20915),
            .I(\PWMInstance6.periodCounterZ0Z_16 ));
    Odrv4 I__3388 (
            .O(N__20912),
            .I(\PWMInstance6.periodCounterZ0Z_16 ));
    InMux I__3387 (
            .O(N__20907),
            .I(N__20904));
    LocalMux I__3386 (
            .O(N__20904),
            .I(data_receivedZ0Z_18));
    InMux I__3385 (
            .O(N__20901),
            .I(N__20898));
    LocalMux I__3384 (
            .O(N__20898),
            .I(data_receivedZ0Z_17));
    InMux I__3383 (
            .O(N__20895),
            .I(N__20892));
    LocalMux I__3382 (
            .O(N__20892),
            .I(data_receivedZ0Z_16));
    InMux I__3381 (
            .O(N__20889),
            .I(N__20885));
    InMux I__3380 (
            .O(N__20888),
            .I(N__20882));
    LocalMux I__3379 (
            .O(N__20885),
            .I(data_receivedZ0Z_15));
    LocalMux I__3378 (
            .O(N__20882),
            .I(data_receivedZ0Z_15));
    InMux I__3377 (
            .O(N__20877),
            .I(N__20872));
    InMux I__3376 (
            .O(N__20876),
            .I(N__20869));
    InMux I__3375 (
            .O(N__20875),
            .I(N__20866));
    LocalMux I__3374 (
            .O(N__20872),
            .I(N__20863));
    LocalMux I__3373 (
            .O(N__20869),
            .I(N__20860));
    LocalMux I__3372 (
            .O(N__20866),
            .I(N__20857));
    Span4Mux_h I__3371 (
            .O(N__20863),
            .I(N__20852));
    Span4Mux_h I__3370 (
            .O(N__20860),
            .I(N__20852));
    Span4Mux_v I__3369 (
            .O(N__20857),
            .I(N__20849));
    Odrv4 I__3368 (
            .O(N__20852),
            .I(dataRead7_11));
    Odrv4 I__3367 (
            .O(N__20849),
            .I(dataRead7_11));
    CascadeMux I__3366 (
            .O(N__20844),
            .I(N__20841));
    InMux I__3365 (
            .O(N__20841),
            .I(N__20837));
    InMux I__3364 (
            .O(N__20840),
            .I(N__20834));
    LocalMux I__3363 (
            .O(N__20837),
            .I(N__20831));
    LocalMux I__3362 (
            .O(N__20834),
            .I(N__20825));
    Span4Mux_v I__3361 (
            .O(N__20831),
            .I(N__20825));
    InMux I__3360 (
            .O(N__20830),
            .I(N__20822));
    Odrv4 I__3359 (
            .O(N__20825),
            .I(dataRead6_11));
    LocalMux I__3358 (
            .O(N__20822),
            .I(dataRead6_11));
    CascadeMux I__3357 (
            .O(N__20817),
            .I(OutReg_ess_RNO_1Z0Z_11_cascade_));
    InMux I__3356 (
            .O(N__20814),
            .I(N__20811));
    LocalMux I__3355 (
            .O(N__20811),
            .I(OutReg_ess_RNO_2Z0Z_11));
    CascadeMux I__3354 (
            .O(N__20808),
            .I(OutReg_ess_RNO_0Z0Z_11_cascade_));
    InMux I__3353 (
            .O(N__20805),
            .I(N__20802));
    LocalMux I__3352 (
            .O(N__20802),
            .I(OutReg_ess_RNO_0Z0Z_13));
    CascadeMux I__3351 (
            .O(N__20799),
            .I(N__20796));
    InMux I__3350 (
            .O(N__20796),
            .I(N__20793));
    LocalMux I__3349 (
            .O(N__20793),
            .I(N__20790));
    Odrv4 I__3348 (
            .O(N__20790),
            .I(\QuadInstance6.Quad_RNI79A91Z0Z_8 ));
    CascadeMux I__3347 (
            .O(N__20787),
            .I(\QuadInstance6.un1_count_enable_i_a2_0_1_cascade_ ));
    CascadeMux I__3346 (
            .O(N__20784),
            .I(N__20781));
    InMux I__3345 (
            .O(N__20781),
            .I(N__20778));
    LocalMux I__3344 (
            .O(N__20778),
            .I(N__20775));
    Odrv12 I__3343 (
            .O(N__20775),
            .I(\QuadInstance6.Quad_RNI35A91Z0Z_4 ));
    CascadeMux I__3342 (
            .O(N__20772),
            .I(N__20769));
    InMux I__3341 (
            .O(N__20769),
            .I(N__20766));
    LocalMux I__3340 (
            .O(N__20766),
            .I(N__20763));
    Odrv4 I__3339 (
            .O(N__20763),
            .I(\QuadInstance6.Quad_RNIIGNB1Z0Z_12 ));
    CascadeMux I__3338 (
            .O(N__20760),
            .I(N__20757));
    InMux I__3337 (
            .O(N__20757),
            .I(N__20754));
    LocalMux I__3336 (
            .O(N__20754),
            .I(N__20751));
    Odrv12 I__3335 (
            .O(N__20751),
            .I(\QuadInstance6.Quad_RNI57A91Z0Z_6 ));
    CascadeMux I__3334 (
            .O(N__20748),
            .I(N__20745));
    InMux I__3333 (
            .O(N__20745),
            .I(N__20742));
    LocalMux I__3332 (
            .O(N__20742),
            .I(N__20739));
    Odrv12 I__3331 (
            .O(N__20739),
            .I(\QuadInstance6.Quad_RNI68A91Z0Z_7 ));
    InMux I__3330 (
            .O(N__20736),
            .I(N__20733));
    LocalMux I__3329 (
            .O(N__20733),
            .I(OutReg_0_4_i_m3_ns_1_13));
    InMux I__3328 (
            .O(N__20730),
            .I(N__20727));
    LocalMux I__3327 (
            .O(N__20727),
            .I(OutReg_ess_RNO_1Z0Z_13));
    InMux I__3326 (
            .O(N__20724),
            .I(N__20721));
    LocalMux I__3325 (
            .O(N__20721),
            .I(N__20718));
    Span4Mux_v I__3324 (
            .O(N__20718),
            .I(N__20715));
    Odrv4 I__3323 (
            .O(N__20715),
            .I(\QuadInstance7.Quad_RNO_0_7_10 ));
    InMux I__3322 (
            .O(N__20712),
            .I(N__20709));
    LocalMux I__3321 (
            .O(N__20709),
            .I(N__20706));
    Odrv4 I__3320 (
            .O(N__20706),
            .I(\QuadInstance5.Quad_RNO_0_5_9 ));
    CascadeMux I__3319 (
            .O(N__20703),
            .I(N__20700));
    InMux I__3318 (
            .O(N__20700),
            .I(N__20697));
    LocalMux I__3317 (
            .O(N__20697),
            .I(N__20694));
    Odrv4 I__3316 (
            .O(N__20694),
            .I(\QuadInstance6.Quad_RNI02A91Z0Z_1 ));
    CascadeMux I__3315 (
            .O(N__20691),
            .I(\QuadInstance6.count_enable_cascade_ ));
    CascadeMux I__3314 (
            .O(N__20688),
            .I(N__20685));
    InMux I__3313 (
            .O(N__20685),
            .I(N__20682));
    LocalMux I__3312 (
            .O(N__20682),
            .I(N__20679));
    Odrv4 I__3311 (
            .O(N__20679),
            .I(\QuadInstance6.Quad_RNI13A91Z0Z_2 ));
    CascadeMux I__3310 (
            .O(N__20676),
            .I(N__20673));
    InMux I__3309 (
            .O(N__20673),
            .I(N__20670));
    LocalMux I__3308 (
            .O(N__20670),
            .I(N__20667));
    Odrv4 I__3307 (
            .O(N__20667),
            .I(\QuadInstance6.Quad_RNIHFNB1Z0Z_11 ));
    CascadeMux I__3306 (
            .O(N__20664),
            .I(N__20661));
    InMux I__3305 (
            .O(N__20661),
            .I(N__20658));
    LocalMux I__3304 (
            .O(N__20658),
            .I(N__20655));
    Odrv4 I__3303 (
            .O(N__20655),
            .I(\QuadInstance6.Quad_RNI24A91Z0Z_3 ));
    CascadeMux I__3302 (
            .O(N__20652),
            .I(N__20649));
    InMux I__3301 (
            .O(N__20649),
            .I(N__20646));
    LocalMux I__3300 (
            .O(N__20646),
            .I(N__20643));
    Odrv4 I__3299 (
            .O(N__20643),
            .I(\QuadInstance6.Quad_RNI46A91Z0Z_5 ));
    CascadeMux I__3298 (
            .O(N__20640),
            .I(N__20637));
    InMux I__3297 (
            .O(N__20637),
            .I(N__20634));
    LocalMux I__3296 (
            .O(N__20634),
            .I(N__20631));
    Odrv4 I__3295 (
            .O(N__20631),
            .I(\QuadInstance6.Quad_RNI8AA91Z0Z_9 ));
    InMux I__3294 (
            .O(N__20628),
            .I(\QuadInstance6.un1_Quad_cry_11 ));
    InMux I__3293 (
            .O(N__20625),
            .I(N__20622));
    LocalMux I__3292 (
            .O(N__20622),
            .I(N__20619));
    Odrv4 I__3291 (
            .O(N__20619),
            .I(\QuadInstance6.Quad_RNO_0_6_13 ));
    InMux I__3290 (
            .O(N__20616),
            .I(\QuadInstance6.un1_Quad_cry_12 ));
    InMux I__3289 (
            .O(N__20613),
            .I(N__20610));
    LocalMux I__3288 (
            .O(N__20610),
            .I(N__20607));
    Odrv12 I__3287 (
            .O(N__20607),
            .I(\QuadInstance6.Quad_RNIKINB1Z0Z_14 ));
    InMux I__3286 (
            .O(N__20604),
            .I(\QuadInstance6.un1_Quad_cry_13 ));
    InMux I__3285 (
            .O(N__20601),
            .I(N__20598));
    LocalMux I__3284 (
            .O(N__20598),
            .I(N__20595));
    Odrv4 I__3283 (
            .O(N__20595),
            .I(\QuadInstance6.un1_Quad_axb_15 ));
    InMux I__3282 (
            .O(N__20592),
            .I(\QuadInstance6.un1_Quad_cry_14 ));
    InMux I__3281 (
            .O(N__20589),
            .I(N__20586));
    LocalMux I__3280 (
            .O(N__20586),
            .I(N__20583));
    Odrv4 I__3279 (
            .O(N__20583),
            .I(\QuadInstance6.Quad_RNO_0_5_1 ));
    InMux I__3278 (
            .O(N__20580),
            .I(N__20577));
    LocalMux I__3277 (
            .O(N__20577),
            .I(N__20574));
    Span4Mux_h I__3276 (
            .O(N__20574),
            .I(N__20571));
    Odrv4 I__3275 (
            .O(N__20571),
            .I(\QuadInstance7.Quad_RNO_0_7_8 ));
    InMux I__3274 (
            .O(N__20568),
            .I(N__20565));
    LocalMux I__3273 (
            .O(N__20565),
            .I(\QuadInstance6.Quad_RNO_0_6_14 ));
    CascadeMux I__3272 (
            .O(N__20562),
            .I(N__20559));
    InMux I__3271 (
            .O(N__20559),
            .I(N__20555));
    InMux I__3270 (
            .O(N__20558),
            .I(N__20551));
    LocalMux I__3269 (
            .O(N__20555),
            .I(N__20548));
    CascadeMux I__3268 (
            .O(N__20554),
            .I(N__20545));
    LocalMux I__3267 (
            .O(N__20551),
            .I(N__20542));
    Span12Mux_s5_v I__3266 (
            .O(N__20548),
            .I(N__20539));
    InMux I__3265 (
            .O(N__20545),
            .I(N__20536));
    Span4Mux_h I__3264 (
            .O(N__20542),
            .I(N__20533));
    Odrv12 I__3263 (
            .O(N__20539),
            .I(dataRead6_14));
    LocalMux I__3262 (
            .O(N__20536),
            .I(dataRead6_14));
    Odrv4 I__3261 (
            .O(N__20533),
            .I(dataRead6_14));
    InMux I__3260 (
            .O(N__20526),
            .I(N__20523));
    LocalMux I__3259 (
            .O(N__20523),
            .I(\QuadInstance6.Quad_RNO_0_6_10 ));
    InMux I__3258 (
            .O(N__20520),
            .I(\QuadInstance6.un1_Quad_cry_3 ));
    InMux I__3257 (
            .O(N__20517),
            .I(N__20514));
    LocalMux I__3256 (
            .O(N__20514),
            .I(\QuadInstance6.Quad_RNO_0_6_5 ));
    InMux I__3255 (
            .O(N__20511),
            .I(\QuadInstance6.un1_Quad_cry_4 ));
    InMux I__3254 (
            .O(N__20508),
            .I(N__20505));
    LocalMux I__3253 (
            .O(N__20505),
            .I(\QuadInstance6.Quad_RNO_0_6_6 ));
    InMux I__3252 (
            .O(N__20502),
            .I(\QuadInstance6.un1_Quad_cry_5 ));
    InMux I__3251 (
            .O(N__20499),
            .I(N__20496));
    LocalMux I__3250 (
            .O(N__20496),
            .I(\QuadInstance6.Quad_RNO_0_6_7 ));
    InMux I__3249 (
            .O(N__20493),
            .I(\QuadInstance6.un1_Quad_cry_6 ));
    InMux I__3248 (
            .O(N__20490),
            .I(N__20487));
    LocalMux I__3247 (
            .O(N__20487),
            .I(\QuadInstance6.Quad_RNO_0_6_8 ));
    InMux I__3246 (
            .O(N__20484),
            .I(bfn_12_6_0_));
    InMux I__3245 (
            .O(N__20481),
            .I(\QuadInstance6.un1_Quad_cry_8 ));
    InMux I__3244 (
            .O(N__20478),
            .I(\QuadInstance6.un1_Quad_cry_9 ));
    InMux I__3243 (
            .O(N__20475),
            .I(N__20472));
    LocalMux I__3242 (
            .O(N__20472),
            .I(\QuadInstance6.Quad_RNO_0_6_11 ));
    InMux I__3241 (
            .O(N__20469),
            .I(\QuadInstance6.un1_Quad_cry_10 ));
    InMux I__3240 (
            .O(N__20466),
            .I(N__20463));
    LocalMux I__3239 (
            .O(N__20463),
            .I(N__20460));
    Odrv4 I__3238 (
            .O(N__20460),
            .I(\QuadInstance6.Quad_RNO_0_6_12 ));
    InMux I__3237 (
            .O(N__20457),
            .I(N__20454));
    LocalMux I__3236 (
            .O(N__20454),
            .I(N__20451));
    Span4Mux_h I__3235 (
            .O(N__20451),
            .I(N__20448));
    Odrv4 I__3234 (
            .O(N__20448),
            .I(\QuadInstance5.Quad_RNO_0_5_5 ));
    InMux I__3233 (
            .O(N__20445),
            .I(N__20442));
    LocalMux I__3232 (
            .O(N__20442),
            .I(N__20439));
    Span4Mux_h I__3231 (
            .O(N__20439),
            .I(N__20436));
    Odrv4 I__3230 (
            .O(N__20436),
            .I(\QuadInstance7.Quad_RNO_0_7_5 ));
    InMux I__3229 (
            .O(N__20433),
            .I(\QuadInstance6.un1_Quad_cry_0 ));
    InMux I__3228 (
            .O(N__20430),
            .I(N__20427));
    LocalMux I__3227 (
            .O(N__20427),
            .I(\QuadInstance6.Quad_RNO_0_6_2 ));
    InMux I__3226 (
            .O(N__20424),
            .I(\QuadInstance6.un1_Quad_cry_1 ));
    InMux I__3225 (
            .O(N__20421),
            .I(N__20418));
    LocalMux I__3224 (
            .O(N__20418),
            .I(\QuadInstance6.Quad_RNO_0_6_3 ));
    InMux I__3223 (
            .O(N__20415),
            .I(\QuadInstance6.un1_Quad_cry_2 ));
    InMux I__3222 (
            .O(N__20412),
            .I(\PWMInstance6.un1_periodCounter_2_cry_12 ));
    InMux I__3221 (
            .O(N__20409),
            .I(\PWMInstance6.un1_periodCounter_2_cry_13 ));
    InMux I__3220 (
            .O(N__20406),
            .I(\PWMInstance6.un1_periodCounter_2_cry_14 ));
    InMux I__3219 (
            .O(N__20403),
            .I(bfn_11_16_0_));
    InMux I__3218 (
            .O(N__20400),
            .I(N__20397));
    LocalMux I__3217 (
            .O(N__20397),
            .I(N__20394));
    Span4Mux_h I__3216 (
            .O(N__20394),
            .I(N__20391));
    Odrv4 I__3215 (
            .O(N__20391),
            .I(ch3_A_c));
    InMux I__3214 (
            .O(N__20388),
            .I(N__20385));
    LocalMux I__3213 (
            .O(N__20385),
            .I(N__20382));
    Span4Mux_v I__3212 (
            .O(N__20382),
            .I(N__20379));
    Span4Mux_v I__3211 (
            .O(N__20379),
            .I(N__20376));
    Span4Mux_v I__3210 (
            .O(N__20376),
            .I(N__20373));
    Odrv4 I__3209 (
            .O(N__20373),
            .I(\QuadInstance3.delayedCh_AZ0Z_0 ));
    InMux I__3208 (
            .O(N__20370),
            .I(N__20367));
    LocalMux I__3207 (
            .O(N__20367),
            .I(N__20364));
    Span4Mux_h I__3206 (
            .O(N__20364),
            .I(N__20361));
    Span4Mux_h I__3205 (
            .O(N__20361),
            .I(N__20358));
    Odrv4 I__3204 (
            .O(N__20358),
            .I(\QuadInstance2.Quad_RNO_0_2_5 ));
    InMux I__3203 (
            .O(N__20355),
            .I(N__20352));
    LocalMux I__3202 (
            .O(N__20352),
            .I(N__20347));
    InMux I__3201 (
            .O(N__20351),
            .I(N__20344));
    InMux I__3200 (
            .O(N__20350),
            .I(N__20341));
    Span4Mux_v I__3199 (
            .O(N__20347),
            .I(N__20338));
    LocalMux I__3198 (
            .O(N__20344),
            .I(\PWMInstance6.periodCounterZ0Z_4 ));
    LocalMux I__3197 (
            .O(N__20341),
            .I(\PWMInstance6.periodCounterZ0Z_4 ));
    Odrv4 I__3196 (
            .O(N__20338),
            .I(\PWMInstance6.periodCounterZ0Z_4 ));
    InMux I__3195 (
            .O(N__20331),
            .I(\PWMInstance6.un1_periodCounter_2_cry_3 ));
    InMux I__3194 (
            .O(N__20328),
            .I(N__20324));
    InMux I__3193 (
            .O(N__20327),
            .I(N__20320));
    LocalMux I__3192 (
            .O(N__20324),
            .I(N__20317));
    InMux I__3191 (
            .O(N__20323),
            .I(N__20314));
    LocalMux I__3190 (
            .O(N__20320),
            .I(\PWMInstance6.periodCounterZ0Z_5 ));
    Odrv4 I__3189 (
            .O(N__20317),
            .I(\PWMInstance6.periodCounterZ0Z_5 ));
    LocalMux I__3188 (
            .O(N__20314),
            .I(\PWMInstance6.periodCounterZ0Z_5 ));
    InMux I__3187 (
            .O(N__20307),
            .I(\PWMInstance6.un1_periodCounter_2_cry_4 ));
    InMux I__3186 (
            .O(N__20304),
            .I(\PWMInstance6.un1_periodCounter_2_cry_5 ));
    InMux I__3185 (
            .O(N__20301),
            .I(\PWMInstance6.un1_periodCounter_2_cry_6 ));
    InMux I__3184 (
            .O(N__20298),
            .I(bfn_11_15_0_));
    InMux I__3183 (
            .O(N__20295),
            .I(\PWMInstance6.un1_periodCounter_2_cry_8 ));
    InMux I__3182 (
            .O(N__20292),
            .I(\PWMInstance6.un1_periodCounter_2_cry_9 ));
    InMux I__3181 (
            .O(N__20289),
            .I(\PWMInstance6.un1_periodCounter_2_cry_10 ));
    InMux I__3180 (
            .O(N__20286),
            .I(\PWMInstance6.un1_periodCounter_2_cry_11 ));
    CascadeMux I__3179 (
            .O(N__20283),
            .I(N__20279));
    CascadeMux I__3178 (
            .O(N__20282),
            .I(N__20276));
    InMux I__3177 (
            .O(N__20279),
            .I(N__20273));
    InMux I__3176 (
            .O(N__20276),
            .I(N__20270));
    LocalMux I__3175 (
            .O(N__20273),
            .I(N__20267));
    LocalMux I__3174 (
            .O(N__20270),
            .I(N__20264));
    Span4Mux_v I__3173 (
            .O(N__20267),
            .I(N__20260));
    Span4Mux_h I__3172 (
            .O(N__20264),
            .I(N__20257));
    InMux I__3171 (
            .O(N__20263),
            .I(N__20254));
    Odrv4 I__3170 (
            .O(N__20260),
            .I(dataRead7_14));
    Odrv4 I__3169 (
            .O(N__20257),
            .I(dataRead7_14));
    LocalMux I__3168 (
            .O(N__20254),
            .I(dataRead7_14));
    CascadeMux I__3167 (
            .O(N__20247),
            .I(OutReg_0_4_i_m3_ns_1_14_cascade_));
    CascadeMux I__3166 (
            .O(N__20244),
            .I(N__20241));
    InMux I__3165 (
            .O(N__20241),
            .I(N__20235));
    InMux I__3164 (
            .O(N__20240),
            .I(N__20235));
    LocalMux I__3163 (
            .O(N__20235),
            .I(pwmWrite_fastZ0Z_5));
    CascadeMux I__3162 (
            .O(N__20232),
            .I(N__20228));
    CascadeMux I__3161 (
            .O(N__20231),
            .I(N__20225));
    InMux I__3160 (
            .O(N__20228),
            .I(N__20217));
    InMux I__3159 (
            .O(N__20225),
            .I(N__20217));
    InMux I__3158 (
            .O(N__20224),
            .I(N__20217));
    LocalMux I__3157 (
            .O(N__20217),
            .I(pwmWriteZ0Z_5));
    InMux I__3156 (
            .O(N__20214),
            .I(\PWMInstance6.un1_periodCounter_2_cry_0 ));
    InMux I__3155 (
            .O(N__20211),
            .I(N__20206));
    InMux I__3154 (
            .O(N__20210),
            .I(N__20203));
    InMux I__3153 (
            .O(N__20209),
            .I(N__20200));
    LocalMux I__3152 (
            .O(N__20206),
            .I(N__20197));
    LocalMux I__3151 (
            .O(N__20203),
            .I(\PWMInstance6.periodCounterZ0Z_2 ));
    LocalMux I__3150 (
            .O(N__20200),
            .I(\PWMInstance6.periodCounterZ0Z_2 ));
    Odrv4 I__3149 (
            .O(N__20197),
            .I(\PWMInstance6.periodCounterZ0Z_2 ));
    InMux I__3148 (
            .O(N__20190),
            .I(\PWMInstance6.un1_periodCounter_2_cry_1 ));
    CascadeMux I__3147 (
            .O(N__20187),
            .I(N__20184));
    InMux I__3146 (
            .O(N__20184),
            .I(N__20181));
    LocalMux I__3145 (
            .O(N__20181),
            .I(N__20176));
    InMux I__3144 (
            .O(N__20180),
            .I(N__20173));
    InMux I__3143 (
            .O(N__20179),
            .I(N__20170));
    Span4Mux_v I__3142 (
            .O(N__20176),
            .I(N__20167));
    LocalMux I__3141 (
            .O(N__20173),
            .I(\PWMInstance6.periodCounterZ0Z_3 ));
    LocalMux I__3140 (
            .O(N__20170),
            .I(\PWMInstance6.periodCounterZ0Z_3 ));
    Odrv4 I__3139 (
            .O(N__20167),
            .I(\PWMInstance6.periodCounterZ0Z_3 ));
    InMux I__3138 (
            .O(N__20160),
            .I(\PWMInstance6.un1_periodCounter_2_cry_2 ));
    InMux I__3137 (
            .O(N__20157),
            .I(N__20154));
    LocalMux I__3136 (
            .O(N__20154),
            .I(\QuadInstance3.Quad_RNO_0_3_14 ));
    InMux I__3135 (
            .O(N__20151),
            .I(N__20148));
    LocalMux I__3134 (
            .O(N__20148),
            .I(N__20145));
    Odrv4 I__3133 (
            .O(N__20145),
            .I(\QuadInstance5.Quad_RNO_0_5_2 ));
    InMux I__3132 (
            .O(N__20142),
            .I(N__20139));
    LocalMux I__3131 (
            .O(N__20139),
            .I(N__20136));
    Odrv4 I__3130 (
            .O(N__20136),
            .I(\QuadInstance7.Quad_RNO_0_7_14 ));
    InMux I__3129 (
            .O(N__20133),
            .I(N__20130));
    LocalMux I__3128 (
            .O(N__20130),
            .I(\QuadInstance3.Quad_RNO_0_3_10 ));
    InMux I__3127 (
            .O(N__20127),
            .I(N__20124));
    LocalMux I__3126 (
            .O(N__20124),
            .I(\QuadInstance3.Quad_RNO_0_3_11 ));
    InMux I__3125 (
            .O(N__20121),
            .I(N__20118));
    LocalMux I__3124 (
            .O(N__20118),
            .I(N__20115));
    Odrv4 I__3123 (
            .O(N__20115),
            .I(OutReg_ess_RNO_2Z0Z_13));
    InMux I__3122 (
            .O(N__20112),
            .I(N__20109));
    LocalMux I__3121 (
            .O(N__20109),
            .I(N__20105));
    InMux I__3120 (
            .O(N__20108),
            .I(N__20102));
    Span4Mux_h I__3119 (
            .O(N__20105),
            .I(N__20098));
    LocalMux I__3118 (
            .O(N__20102),
            .I(N__20095));
    InMux I__3117 (
            .O(N__20101),
            .I(N__20092));
    Span4Mux_h I__3116 (
            .O(N__20098),
            .I(N__20087));
    Span4Mux_h I__3115 (
            .O(N__20095),
            .I(N__20087));
    LocalMux I__3114 (
            .O(N__20092),
            .I(dataRead5_11));
    Odrv4 I__3113 (
            .O(N__20087),
            .I(dataRead5_11));
    CascadeMux I__3112 (
            .O(N__20082),
            .I(OutReg_0_5_i_m3_i_m3_ns_1_11_cascade_));
    CascadeMux I__3111 (
            .O(N__20079),
            .I(N__20076));
    InMux I__3110 (
            .O(N__20076),
            .I(N__20073));
    LocalMux I__3109 (
            .O(N__20073),
            .I(N__20069));
    CascadeMux I__3108 (
            .O(N__20072),
            .I(N__20066));
    Span4Mux_v I__3107 (
            .O(N__20069),
            .I(N__20062));
    InMux I__3106 (
            .O(N__20066),
            .I(N__20059));
    InMux I__3105 (
            .O(N__20065),
            .I(N__20056));
    Odrv4 I__3104 (
            .O(N__20062),
            .I(dataRead3_14));
    LocalMux I__3103 (
            .O(N__20059),
            .I(dataRead3_14));
    LocalMux I__3102 (
            .O(N__20056),
            .I(dataRead3_14));
    CascadeMux I__3101 (
            .O(N__20049),
            .I(N__20044));
    InMux I__3100 (
            .O(N__20048),
            .I(N__20041));
    CascadeMux I__3099 (
            .O(N__20047),
            .I(N__20038));
    InMux I__3098 (
            .O(N__20044),
            .I(N__20035));
    LocalMux I__3097 (
            .O(N__20041),
            .I(N__20032));
    InMux I__3096 (
            .O(N__20038),
            .I(N__20029));
    LocalMux I__3095 (
            .O(N__20035),
            .I(N__20024));
    Span4Mux_h I__3094 (
            .O(N__20032),
            .I(N__20024));
    LocalMux I__3093 (
            .O(N__20029),
            .I(dataRead2_14));
    Odrv4 I__3092 (
            .O(N__20024),
            .I(dataRead2_14));
    CascadeMux I__3091 (
            .O(N__20019),
            .I(N__20016));
    InMux I__3090 (
            .O(N__20016),
            .I(N__20013));
    LocalMux I__3089 (
            .O(N__20013),
            .I(N__20009));
    CascadeMux I__3088 (
            .O(N__20012),
            .I(N__20005));
    Span4Mux_v I__3087 (
            .O(N__20009),
            .I(N__20002));
    InMux I__3086 (
            .O(N__20008),
            .I(N__19999));
    InMux I__3085 (
            .O(N__20005),
            .I(N__19996));
    Span4Mux_h I__3084 (
            .O(N__20002),
            .I(N__19993));
    LocalMux I__3083 (
            .O(N__19999),
            .I(dataRead5_13));
    LocalMux I__3082 (
            .O(N__19996),
            .I(dataRead5_13));
    Odrv4 I__3081 (
            .O(N__19993),
            .I(dataRead5_13));
    InMux I__3080 (
            .O(N__19986),
            .I(N__19983));
    LocalMux I__3079 (
            .O(N__19983),
            .I(N__19980));
    Span4Mux_v I__3078 (
            .O(N__19980),
            .I(N__19977));
    Odrv4 I__3077 (
            .O(N__19977),
            .I(\QuadInstance2.Quad_RNO_0_2_13 ));
    InMux I__3076 (
            .O(N__19974),
            .I(N__19970));
    InMux I__3075 (
            .O(N__19973),
            .I(N__19967));
    LocalMux I__3074 (
            .O(N__19970),
            .I(N__19964));
    LocalMux I__3073 (
            .O(N__19967),
            .I(N__19961));
    Span4Mux_v I__3072 (
            .O(N__19964),
            .I(N__19957));
    Span4Mux_h I__3071 (
            .O(N__19961),
            .I(N__19954));
    InMux I__3070 (
            .O(N__19960),
            .I(N__19951));
    Odrv4 I__3069 (
            .O(N__19957),
            .I(dataRead2_13));
    Odrv4 I__3068 (
            .O(N__19954),
            .I(dataRead2_13));
    LocalMux I__3067 (
            .O(N__19951),
            .I(dataRead2_13));
    InMux I__3066 (
            .O(N__19944),
            .I(N__19941));
    LocalMux I__3065 (
            .O(N__19941),
            .I(\QuadInstance3.Quad_RNO_0_3_13 ));
    CascadeMux I__3064 (
            .O(N__19938),
            .I(N__19935));
    InMux I__3063 (
            .O(N__19935),
            .I(N__19932));
    LocalMux I__3062 (
            .O(N__19932),
            .I(N__19929));
    Span4Mux_v I__3061 (
            .O(N__19929),
            .I(N__19925));
    InMux I__3060 (
            .O(N__19928),
            .I(N__19922));
    Sp12to4 I__3059 (
            .O(N__19925),
            .I(N__19918));
    LocalMux I__3058 (
            .O(N__19922),
            .I(N__19915));
    InMux I__3057 (
            .O(N__19921),
            .I(N__19912));
    Odrv12 I__3056 (
            .O(N__19918),
            .I(dataRead3_13));
    Odrv4 I__3055 (
            .O(N__19915),
            .I(dataRead3_13));
    LocalMux I__3054 (
            .O(N__19912),
            .I(dataRead3_13));
    InMux I__3053 (
            .O(N__19905),
            .I(N__19902));
    LocalMux I__3052 (
            .O(N__19902),
            .I(\QuadInstance3.Quad_RNO_0_3_12 ));
    CascadeMux I__3051 (
            .O(N__19899),
            .I(N__19896));
    InMux I__3050 (
            .O(N__19896),
            .I(N__19893));
    LocalMux I__3049 (
            .O(N__19893),
            .I(\QuadInstance3.Quad_RNO_0_3_8 ));
    InMux I__3048 (
            .O(N__19890),
            .I(N__19887));
    LocalMux I__3047 (
            .O(N__19887),
            .I(N__19884));
    Span4Mux_h I__3046 (
            .O(N__19884),
            .I(N__19881));
    Odrv4 I__3045 (
            .O(N__19881),
            .I(\QuadInstance7.Quad_RNO_0_7_7 ));
    InMux I__3044 (
            .O(N__19878),
            .I(N__19875));
    LocalMux I__3043 (
            .O(N__19875),
            .I(N__19872));
    Odrv12 I__3042 (
            .O(N__19872),
            .I(\QuadInstance2.Quad_RNO_0_2_11 ));
    InMux I__3041 (
            .O(N__19869),
            .I(N__19866));
    LocalMux I__3040 (
            .O(N__19866),
            .I(\QuadInstance5.Quad_RNO_0_5_10 ));
    InMux I__3039 (
            .O(N__19863),
            .I(N__19860));
    LocalMux I__3038 (
            .O(N__19860),
            .I(\QuadInstance5.Quad_RNO_0_5_11 ));
    InMux I__3037 (
            .O(N__19857),
            .I(N__19854));
    LocalMux I__3036 (
            .O(N__19854),
            .I(N__19851));
    Span4Mux_h I__3035 (
            .O(N__19851),
            .I(N__19848));
    Odrv4 I__3034 (
            .O(N__19848),
            .I(\QuadInstance2.Quad_RNO_0_2_8 ));
    InMux I__3033 (
            .O(N__19845),
            .I(N__19842));
    LocalMux I__3032 (
            .O(N__19842),
            .I(N__19839));
    Odrv4 I__3031 (
            .O(N__19839),
            .I(\QuadInstance3.Quad_RNO_0_3_9 ));
    InMux I__3030 (
            .O(N__19836),
            .I(N__19833));
    LocalMux I__3029 (
            .O(N__19833),
            .I(N__19830));
    Span4Mux_h I__3028 (
            .O(N__19830),
            .I(N__19827));
    Odrv4 I__3027 (
            .O(N__19827),
            .I(\QuadInstance7.Quad_RNO_0_7_9 ));
    InMux I__3026 (
            .O(N__19824),
            .I(N__19821));
    LocalMux I__3025 (
            .O(N__19821),
            .I(N__19818));
    Odrv4 I__3024 (
            .O(N__19818),
            .I(\QuadInstance5.Quad_RNO_0_5_8 ));
    InMux I__3023 (
            .O(N__19815),
            .I(N__19812));
    LocalMux I__3022 (
            .O(N__19812),
            .I(N__19809));
    Span4Mux_v I__3021 (
            .O(N__19809),
            .I(N__19806));
    Odrv4 I__3020 (
            .O(N__19806),
            .I(\QuadInstance3.Quad_RNO_0_3_3 ));
    InMux I__3019 (
            .O(N__19803),
            .I(N__19800));
    LocalMux I__3018 (
            .O(N__19800),
            .I(N__19797));
    Odrv12 I__3017 (
            .O(N__19797),
            .I(\QuadInstance2.Quad_RNO_0_2_7 ));
    InMux I__3016 (
            .O(N__19794),
            .I(N__19791));
    LocalMux I__3015 (
            .O(N__19791),
            .I(N__19788));
    Odrv4 I__3014 (
            .O(N__19788),
            .I(\QuadInstance3.Quad_RNO_0_3_7 ));
    InMux I__3013 (
            .O(N__19785),
            .I(N__19782));
    LocalMux I__3012 (
            .O(N__19782),
            .I(\QuadInstance5.Quad_RNO_0_5_7 ));
    InMux I__3011 (
            .O(N__19779),
            .I(N__19776));
    LocalMux I__3010 (
            .O(N__19776),
            .I(N__19773));
    Odrv4 I__3009 (
            .O(N__19773),
            .I(\QuadInstance3.Quad_RNO_0_3_5 ));
    InMux I__3008 (
            .O(N__19770),
            .I(N__19767));
    LocalMux I__3007 (
            .O(N__19767),
            .I(N__19764));
    Span4Mux_h I__3006 (
            .O(N__19764),
            .I(N__19761));
    Odrv4 I__3005 (
            .O(N__19761),
            .I(\QuadInstance2.Quad_RNO_0_2_6 ));
    InMux I__3004 (
            .O(N__19758),
            .I(N__19755));
    LocalMux I__3003 (
            .O(N__19755),
            .I(N__19752));
    Span4Mux_h I__3002 (
            .O(N__19752),
            .I(N__19749));
    Odrv4 I__3001 (
            .O(N__19749),
            .I(\QuadInstance7.Quad_RNO_0_7_2 ));
    InMux I__3000 (
            .O(N__19746),
            .I(N__19743));
    LocalMux I__2999 (
            .O(N__19743),
            .I(N__19740));
    Span4Mux_v I__2998 (
            .O(N__19740),
            .I(N__19737));
    Odrv4 I__2997 (
            .O(N__19737),
            .I(\QuadInstance2.Quad_RNO_0_2_3 ));
    InMux I__2996 (
            .O(N__19734),
            .I(N__19731));
    LocalMux I__2995 (
            .O(N__19731),
            .I(\QuadInstance5.Quad_RNO_0_5_4 ));
    InMux I__2994 (
            .O(N__19728),
            .I(N__19725));
    LocalMux I__2993 (
            .O(N__19725),
            .I(\QuadInstance5.Quad_RNO_0_5_6 ));
    InMux I__2992 (
            .O(N__19722),
            .I(N__19719));
    LocalMux I__2991 (
            .O(N__19719),
            .I(N__19716));
    Span4Mux_h I__2990 (
            .O(N__19716),
            .I(N__19713));
    Odrv4 I__2989 (
            .O(N__19713),
            .I(\QuadInstance7.Quad_RNO_0_7_6 ));
    CascadeMux I__2988 (
            .O(N__19710),
            .I(\PWMInstance6.un1_periodCounter12_1_0_a2_0_0_cascade_ ));
    CascadeMux I__2987 (
            .O(N__19707),
            .I(\PWMInstance6.un1_periodCounter12_1_0_a2_0_12_cascade_ ));
    InMux I__2986 (
            .O(N__19704),
            .I(N__19701));
    LocalMux I__2985 (
            .O(N__19701),
            .I(\PWMInstance6.un1_periodCounter12_1_0_a2_0_10 ));
    InMux I__2984 (
            .O(N__19698),
            .I(N__19695));
    LocalMux I__2983 (
            .O(N__19695),
            .I(\PWMInstance6.PWMPulseWidthCountZ0Z_2 ));
    InMux I__2982 (
            .O(N__19692),
            .I(N__19689));
    LocalMux I__2981 (
            .O(N__19689),
            .I(\PWMInstance6.PWMPulseWidthCountZ0Z_3 ));
    CascadeMux I__2980 (
            .O(N__19686),
            .I(N__19683));
    InMux I__2979 (
            .O(N__19683),
            .I(N__19680));
    LocalMux I__2978 (
            .O(N__19680),
            .I(\PWMInstance6.PWMPulseWidthCountZ0Z_4 ));
    InMux I__2977 (
            .O(N__19677),
            .I(N__19674));
    LocalMux I__2976 (
            .O(N__19674),
            .I(N__19671));
    Span4Mux_v I__2975 (
            .O(N__19671),
            .I(N__19668));
    Odrv4 I__2974 (
            .O(N__19668),
            .I(\QuadInstance2.Quad_RNO_0_2_2 ));
    InMux I__2973 (
            .O(N__19665),
            .I(N__19662));
    LocalMux I__2972 (
            .O(N__19662),
            .I(N__19659));
    Span4Mux_h I__2971 (
            .O(N__19659),
            .I(N__19656));
    Odrv4 I__2970 (
            .O(N__19656),
            .I(\QuadInstance3.Quad_RNO_0_3_2 ));
    CEMux I__2969 (
            .O(N__19653),
            .I(N__19646));
    CEMux I__2968 (
            .O(N__19652),
            .I(N__19643));
    CEMux I__2967 (
            .O(N__19651),
            .I(N__19640));
    CEMux I__2966 (
            .O(N__19650),
            .I(N__19636));
    CEMux I__2965 (
            .O(N__19649),
            .I(N__19632));
    LocalMux I__2964 (
            .O(N__19646),
            .I(N__19627));
    LocalMux I__2963 (
            .O(N__19643),
            .I(N__19627));
    LocalMux I__2962 (
            .O(N__19640),
            .I(N__19624));
    CEMux I__2961 (
            .O(N__19639),
            .I(N__19621));
    LocalMux I__2960 (
            .O(N__19636),
            .I(N__19618));
    CEMux I__2959 (
            .O(N__19635),
            .I(N__19615));
    LocalMux I__2958 (
            .O(N__19632),
            .I(N__19612));
    Span4Mux_v I__2957 (
            .O(N__19627),
            .I(N__19609));
    Span4Mux_v I__2956 (
            .O(N__19624),
            .I(N__19606));
    LocalMux I__2955 (
            .O(N__19621),
            .I(N__19603));
    Span4Mux_h I__2954 (
            .O(N__19618),
            .I(N__19598));
    LocalMux I__2953 (
            .O(N__19615),
            .I(N__19598));
    Span4Mux_h I__2952 (
            .O(N__19612),
            .I(N__19594));
    Span4Mux_h I__2951 (
            .O(N__19609),
            .I(N__19587));
    Span4Mux_h I__2950 (
            .O(N__19606),
            .I(N__19587));
    Span4Mux_v I__2949 (
            .O(N__19603),
            .I(N__19587));
    Span4Mux_h I__2948 (
            .O(N__19598),
            .I(N__19584));
    CEMux I__2947 (
            .O(N__19597),
            .I(N__19581));
    Odrv4 I__2946 (
            .O(N__19594),
            .I(\PWMInstance5.pwmWrite_0_5 ));
    Odrv4 I__2945 (
            .O(N__19587),
            .I(\PWMInstance5.pwmWrite_0_5 ));
    Odrv4 I__2944 (
            .O(N__19584),
            .I(\PWMInstance5.pwmWrite_0_5 ));
    LocalMux I__2943 (
            .O(N__19581),
            .I(\PWMInstance5.pwmWrite_0_5 ));
    InMux I__2942 (
            .O(N__19572),
            .I(N__19562));
    InMux I__2941 (
            .O(N__19571),
            .I(N__19562));
    InMux I__2940 (
            .O(N__19570),
            .I(N__19562));
    InMux I__2939 (
            .O(N__19569),
            .I(N__19559));
    LocalMux I__2938 (
            .O(N__19562),
            .I(\PWMInstance5.clkCountZ0Z_1 ));
    LocalMux I__2937 (
            .O(N__19559),
            .I(\PWMInstance5.clkCountZ0Z_1 ));
    InMux I__2936 (
            .O(N__19554),
            .I(N__19542));
    InMux I__2935 (
            .O(N__19553),
            .I(N__19542));
    InMux I__2934 (
            .O(N__19552),
            .I(N__19542));
    InMux I__2933 (
            .O(N__19551),
            .I(N__19542));
    LocalMux I__2932 (
            .O(N__19542),
            .I(\PWMInstance5.clkCountZ0Z_0 ));
    CascadeMux I__2931 (
            .O(N__19539),
            .I(N__19535));
    InMux I__2930 (
            .O(N__19538),
            .I(N__19532));
    InMux I__2929 (
            .O(N__19535),
            .I(N__19529));
    LocalMux I__2928 (
            .O(N__19532),
            .I(\PWMInstance5.periodCounter12 ));
    LocalMux I__2927 (
            .O(N__19529),
            .I(\PWMInstance5.periodCounter12 ));
    CascadeMux I__2926 (
            .O(N__19524),
            .I(N__19520));
    InMux I__2925 (
            .O(N__19523),
            .I(N__19516));
    InMux I__2924 (
            .O(N__19520),
            .I(N__19513));
    InMux I__2923 (
            .O(N__19519),
            .I(N__19510));
    LocalMux I__2922 (
            .O(N__19516),
            .I(\PWMInstance5.periodCounterZ0Z_15 ));
    LocalMux I__2921 (
            .O(N__19513),
            .I(\PWMInstance5.periodCounterZ0Z_15 ));
    LocalMux I__2920 (
            .O(N__19510),
            .I(\PWMInstance5.periodCounterZ0Z_15 ));
    CascadeMux I__2919 (
            .O(N__19503),
            .I(N__19498));
    InMux I__2918 (
            .O(N__19502),
            .I(N__19495));
    InMux I__2917 (
            .O(N__19501),
            .I(N__19492));
    InMux I__2916 (
            .O(N__19498),
            .I(N__19489));
    LocalMux I__2915 (
            .O(N__19495),
            .I(\PWMInstance5.periodCounterZ0Z_1 ));
    LocalMux I__2914 (
            .O(N__19492),
            .I(\PWMInstance5.periodCounterZ0Z_1 ));
    LocalMux I__2913 (
            .O(N__19489),
            .I(\PWMInstance5.periodCounterZ0Z_1 ));
    CascadeMux I__2912 (
            .O(N__19482),
            .I(\PWMInstance5.periodCounter12_cascade_ ));
    InMux I__2911 (
            .O(N__19479),
            .I(N__19476));
    LocalMux I__2910 (
            .O(N__19476),
            .I(N__19473));
    Odrv4 I__2909 (
            .O(N__19473),
            .I(\PWMInstance5.un1_periodCounter12_1_0_a2_0_9 ));
    CascadeMux I__2908 (
            .O(N__19470),
            .I(\PWMInstance5.un1_periodCounter12_1_0_a2_0_14_cascade_ ));
    InMux I__2907 (
            .O(N__19467),
            .I(N__19464));
    LocalMux I__2906 (
            .O(N__19464),
            .I(\PWMInstance5.un1_periodCounter12_1_0_a2_0_12 ));
    CascadeMux I__2905 (
            .O(N__19461),
            .I(N__19458));
    InMux I__2904 (
            .O(N__19458),
            .I(N__19455));
    LocalMux I__2903 (
            .O(N__19455),
            .I(N__19447));
    InMux I__2902 (
            .O(N__19454),
            .I(N__19442));
    InMux I__2901 (
            .O(N__19453),
            .I(N__19442));
    InMux I__2900 (
            .O(N__19452),
            .I(N__19439));
    InMux I__2899 (
            .O(N__19451),
            .I(N__19436));
    InMux I__2898 (
            .O(N__19450),
            .I(N__19433));
    Span12Mux_v I__2897 (
            .O(N__19447),
            .I(N__19430));
    LocalMux I__2896 (
            .O(N__19442),
            .I(\PWMInstance5.out_0_sqmuxa ));
    LocalMux I__2895 (
            .O(N__19439),
            .I(\PWMInstance5.out_0_sqmuxa ));
    LocalMux I__2894 (
            .O(N__19436),
            .I(\PWMInstance5.out_0_sqmuxa ));
    LocalMux I__2893 (
            .O(N__19433),
            .I(\PWMInstance5.out_0_sqmuxa ));
    Odrv12 I__2892 (
            .O(N__19430),
            .I(\PWMInstance5.out_0_sqmuxa ));
    CascadeMux I__2891 (
            .O(N__19419),
            .I(N__19416));
    InMux I__2890 (
            .O(N__19416),
            .I(N__19411));
    InMux I__2889 (
            .O(N__19415),
            .I(N__19408));
    InMux I__2888 (
            .O(N__19414),
            .I(N__19405));
    LocalMux I__2887 (
            .O(N__19411),
            .I(N__19402));
    LocalMux I__2886 (
            .O(N__19408),
            .I(\PWMInstance5.periodCounterZ0Z_9 ));
    LocalMux I__2885 (
            .O(N__19405),
            .I(\PWMInstance5.periodCounterZ0Z_9 ));
    Odrv12 I__2884 (
            .O(N__19402),
            .I(\PWMInstance5.periodCounterZ0Z_9 ));
    InMux I__2883 (
            .O(N__19395),
            .I(N__19390));
    CascadeMux I__2882 (
            .O(N__19394),
            .I(N__19387));
    InMux I__2881 (
            .O(N__19393),
            .I(N__19384));
    LocalMux I__2880 (
            .O(N__19390),
            .I(N__19381));
    InMux I__2879 (
            .O(N__19387),
            .I(N__19378));
    LocalMux I__2878 (
            .O(N__19384),
            .I(\PWMInstance5.periodCounterZ0Z_5 ));
    Odrv4 I__2877 (
            .O(N__19381),
            .I(\PWMInstance5.periodCounterZ0Z_5 ));
    LocalMux I__2876 (
            .O(N__19378),
            .I(\PWMInstance5.periodCounterZ0Z_5 ));
    CascadeMux I__2875 (
            .O(N__19371),
            .I(N__19366));
    CascadeMux I__2874 (
            .O(N__19370),
            .I(N__19363));
    InMux I__2873 (
            .O(N__19369),
            .I(N__19360));
    InMux I__2872 (
            .O(N__19366),
            .I(N__19357));
    InMux I__2871 (
            .O(N__19363),
            .I(N__19354));
    LocalMux I__2870 (
            .O(N__19360),
            .I(\PWMInstance5.periodCounterZ0Z_11 ));
    LocalMux I__2869 (
            .O(N__19357),
            .I(\PWMInstance5.periodCounterZ0Z_11 ));
    LocalMux I__2868 (
            .O(N__19354),
            .I(\PWMInstance5.periodCounterZ0Z_11 ));
    InMux I__2867 (
            .O(N__19347),
            .I(N__19342));
    CascadeMux I__2866 (
            .O(N__19346),
            .I(N__19339));
    InMux I__2865 (
            .O(N__19345),
            .I(N__19336));
    LocalMux I__2864 (
            .O(N__19342),
            .I(N__19333));
    InMux I__2863 (
            .O(N__19339),
            .I(N__19330));
    LocalMux I__2862 (
            .O(N__19336),
            .I(\PWMInstance5.periodCounterZ0Z_3 ));
    Odrv4 I__2861 (
            .O(N__19333),
            .I(\PWMInstance5.periodCounterZ0Z_3 ));
    LocalMux I__2860 (
            .O(N__19330),
            .I(\PWMInstance5.periodCounterZ0Z_3 ));
    InMux I__2859 (
            .O(N__19323),
            .I(N__19320));
    LocalMux I__2858 (
            .O(N__19320),
            .I(\PWMInstance5.un1_periodCounter12_1_0_a2_0_10 ));
    InMux I__2857 (
            .O(N__19317),
            .I(N__19312));
    InMux I__2856 (
            .O(N__19316),
            .I(N__19309));
    InMux I__2855 (
            .O(N__19315),
            .I(N__19306));
    LocalMux I__2854 (
            .O(N__19312),
            .I(\PWMInstance5.periodCounterZ0Z_16 ));
    LocalMux I__2853 (
            .O(N__19309),
            .I(\PWMInstance5.periodCounterZ0Z_16 ));
    LocalMux I__2852 (
            .O(N__19306),
            .I(\PWMInstance5.periodCounterZ0Z_16 ));
    InMux I__2851 (
            .O(N__19299),
            .I(N__19294));
    InMux I__2850 (
            .O(N__19298),
            .I(N__19291));
    InMux I__2849 (
            .O(N__19297),
            .I(N__19288));
    LocalMux I__2848 (
            .O(N__19294),
            .I(N__19285));
    LocalMux I__2847 (
            .O(N__19291),
            .I(\PWMInstance5.periodCounterZ0Z_7 ));
    LocalMux I__2846 (
            .O(N__19288),
            .I(\PWMInstance5.periodCounterZ0Z_7 ));
    Odrv4 I__2845 (
            .O(N__19285),
            .I(\PWMInstance5.periodCounterZ0Z_7 ));
    InMux I__2844 (
            .O(N__19278),
            .I(N__19275));
    LocalMux I__2843 (
            .O(N__19275),
            .I(\PWMInstance5.un1_periodCounter12_1_0_a2_0_6 ));
    InMux I__2842 (
            .O(N__19272),
            .I(N__19269));
    LocalMux I__2841 (
            .O(N__19269),
            .I(N__19266));
    Span4Mux_h I__2840 (
            .O(N__19266),
            .I(N__19263));
    Span4Mux_v I__2839 (
            .O(N__19263),
            .I(N__19260));
    Odrv4 I__2838 (
            .O(N__19260),
            .I(\PWMInstance5.un1_PWMPulseWidthCount_0_I_15_c_RNO_4 ));
    InMux I__2837 (
            .O(N__19257),
            .I(N__19252));
    InMux I__2836 (
            .O(N__19256),
            .I(N__19249));
    InMux I__2835 (
            .O(N__19255),
            .I(N__19246));
    LocalMux I__2834 (
            .O(N__19252),
            .I(\PWMInstance5.periodCounterZ0Z_2 ));
    LocalMux I__2833 (
            .O(N__19249),
            .I(\PWMInstance5.periodCounterZ0Z_2 ));
    LocalMux I__2832 (
            .O(N__19246),
            .I(\PWMInstance5.periodCounterZ0Z_2 ));
    InMux I__2831 (
            .O(N__19239),
            .I(N__19234));
    InMux I__2830 (
            .O(N__19238),
            .I(N__19231));
    InMux I__2829 (
            .O(N__19237),
            .I(N__19228));
    LocalMux I__2828 (
            .O(N__19234),
            .I(\PWMInstance5.periodCounterZ0Z_14 ));
    LocalMux I__2827 (
            .O(N__19231),
            .I(\PWMInstance5.periodCounterZ0Z_14 ));
    LocalMux I__2826 (
            .O(N__19228),
            .I(\PWMInstance5.periodCounterZ0Z_14 ));
    InMux I__2825 (
            .O(N__19221),
            .I(N__19216));
    InMux I__2824 (
            .O(N__19220),
            .I(N__19213));
    InMux I__2823 (
            .O(N__19219),
            .I(N__19210));
    LocalMux I__2822 (
            .O(N__19216),
            .I(\PWMInstance5.periodCounterZ0Z_12 ));
    LocalMux I__2821 (
            .O(N__19213),
            .I(\PWMInstance5.periodCounterZ0Z_12 ));
    LocalMux I__2820 (
            .O(N__19210),
            .I(\PWMInstance5.periodCounterZ0Z_12 ));
    CascadeMux I__2819 (
            .O(N__19203),
            .I(\PWMInstance5.un1_periodCounter12_1_0_a2_0_0_cascade_ ));
    InMux I__2818 (
            .O(N__19200),
            .I(N__19195));
    InMux I__2817 (
            .O(N__19199),
            .I(N__19190));
    InMux I__2816 (
            .O(N__19198),
            .I(N__19190));
    LocalMux I__2815 (
            .O(N__19195),
            .I(\PWMInstance5.periodCounterZ0Z_4 ));
    LocalMux I__2814 (
            .O(N__19190),
            .I(\PWMInstance5.periodCounterZ0Z_4 ));
    InMux I__2813 (
            .O(N__19185),
            .I(N__19182));
    LocalMux I__2812 (
            .O(N__19182),
            .I(\PWMInstance5.PWMPulseWidthCountZ0Z_4 ));
    InMux I__2811 (
            .O(N__19179),
            .I(N__19176));
    LocalMux I__2810 (
            .O(N__19176),
            .I(\PWMInstance5.PWMPulseWidthCountZ0Z_5 ));
    InMux I__2809 (
            .O(N__19173),
            .I(N__19168));
    InMux I__2808 (
            .O(N__19172),
            .I(N__19163));
    InMux I__2807 (
            .O(N__19171),
            .I(N__19163));
    LocalMux I__2806 (
            .O(N__19168),
            .I(\PWMInstance5.periodCounterZ0Z_10 ));
    LocalMux I__2805 (
            .O(N__19163),
            .I(\PWMInstance5.periodCounterZ0Z_10 ));
    InMux I__2804 (
            .O(N__19158),
            .I(N__19155));
    LocalMux I__2803 (
            .O(N__19155),
            .I(N__19152));
    Span4Mux_h I__2802 (
            .O(N__19152),
            .I(N__19149));
    Span4Mux_h I__2801 (
            .O(N__19149),
            .I(N__19146));
    Odrv4 I__2800 (
            .O(N__19146),
            .I(\PWMInstance5.PWMPulseWidthCountZ0Z_10 ));
    InMux I__2799 (
            .O(N__19143),
            .I(N__19140));
    LocalMux I__2798 (
            .O(N__19140),
            .I(N__19137));
    Span4Mux_h I__2797 (
            .O(N__19137),
            .I(N__19134));
    Span4Mux_v I__2796 (
            .O(N__19134),
            .I(N__19131));
    Odrv4 I__2795 (
            .O(N__19131),
            .I(\PWMInstance5.un1_PWMPulseWidthCount_0_I_33_c_RNO_4 ));
    InMux I__2794 (
            .O(N__19128),
            .I(N__19125));
    LocalMux I__2793 (
            .O(N__19125),
            .I(\PWMInstance5.PWMPulseWidthCountZ0Z_11 ));
    InMux I__2792 (
            .O(N__19122),
            .I(N__19119));
    LocalMux I__2791 (
            .O(N__19119),
            .I(N__19116));
    Span4Mux_h I__2790 (
            .O(N__19116),
            .I(N__19113));
    Span4Mux_v I__2789 (
            .O(N__19113),
            .I(N__19110));
    Odrv4 I__2788 (
            .O(N__19110),
            .I(\PWMInstance5.un1_periodCounter12_1_0_a2_0 ));
    InMux I__2787 (
            .O(N__19107),
            .I(N__19104));
    LocalMux I__2786 (
            .O(N__19104),
            .I(N__19101));
    Odrv4 I__2785 (
            .O(N__19101),
            .I(\QuadInstance3.Quad_RNIBRAL1Z0Z_4 ));
    InMux I__2784 (
            .O(N__19098),
            .I(N__19095));
    LocalMux I__2783 (
            .O(N__19095),
            .I(N__19092));
    Odrv4 I__2782 (
            .O(N__19092),
            .I(\QuadInstance3.Quad_RNIS50J1Z0Z_14 ));
    CascadeMux I__2781 (
            .O(N__19089),
            .I(N__19085));
    CascadeMux I__2780 (
            .O(N__19088),
            .I(N__19082));
    InMux I__2779 (
            .O(N__19085),
            .I(N__19077));
    InMux I__2778 (
            .O(N__19082),
            .I(N__19077));
    LocalMux I__2777 (
            .O(N__19077),
            .I(\QuadInstance3.delayedCh_BZ0Z_2 ));
    InMux I__2776 (
            .O(N__19074),
            .I(N__19071));
    LocalMux I__2775 (
            .O(N__19071),
            .I(\QuadInstance3.delayedCh_AZ0Z_2 ));
    InMux I__2774 (
            .O(N__19068),
            .I(N__19063));
    InMux I__2773 (
            .O(N__19067),
            .I(N__19058));
    InMux I__2772 (
            .O(N__19066),
            .I(N__19058));
    LocalMux I__2771 (
            .O(N__19063),
            .I(\QuadInstance3.delayedCh_AZ0Z_1 ));
    LocalMux I__2770 (
            .O(N__19058),
            .I(\QuadInstance3.delayedCh_AZ0Z_1 ));
    CascadeMux I__2769 (
            .O(N__19053),
            .I(N__19050));
    InMux I__2768 (
            .O(N__19050),
            .I(N__19047));
    LocalMux I__2767 (
            .O(N__19047),
            .I(N__19044));
    Odrv4 I__2766 (
            .O(N__19044),
            .I(\QuadInstance3.Quad_RNIEUAL1Z0Z_7 ));
    CascadeMux I__2765 (
            .O(N__19041),
            .I(N__19036));
    CascadeMux I__2764 (
            .O(N__19040),
            .I(N__19031));
    InMux I__2763 (
            .O(N__19039),
            .I(N__19015));
    InMux I__2762 (
            .O(N__19036),
            .I(N__19015));
    InMux I__2761 (
            .O(N__19035),
            .I(N__19015));
    InMux I__2760 (
            .O(N__19034),
            .I(N__19008));
    InMux I__2759 (
            .O(N__19031),
            .I(N__19008));
    InMux I__2758 (
            .O(N__19030),
            .I(N__19008));
    InMux I__2757 (
            .O(N__19029),
            .I(N__19001));
    InMux I__2756 (
            .O(N__19028),
            .I(N__19001));
    InMux I__2755 (
            .O(N__19027),
            .I(N__19001));
    InMux I__2754 (
            .O(N__19026),
            .I(N__18994));
    InMux I__2753 (
            .O(N__19025),
            .I(N__18994));
    InMux I__2752 (
            .O(N__19024),
            .I(N__18994));
    InMux I__2751 (
            .O(N__19023),
            .I(N__18989));
    InMux I__2750 (
            .O(N__19022),
            .I(N__18989));
    LocalMux I__2749 (
            .O(N__19015),
            .I(\QuadInstance3.un1_count_enable_i_a2_0_1 ));
    LocalMux I__2748 (
            .O(N__19008),
            .I(\QuadInstance3.un1_count_enable_i_a2_0_1 ));
    LocalMux I__2747 (
            .O(N__19001),
            .I(\QuadInstance3.un1_count_enable_i_a2_0_1 ));
    LocalMux I__2746 (
            .O(N__18994),
            .I(\QuadInstance3.un1_count_enable_i_a2_0_1 ));
    LocalMux I__2745 (
            .O(N__18989),
            .I(\QuadInstance3.un1_count_enable_i_a2_0_1 ));
    InMux I__2744 (
            .O(N__18978),
            .I(N__18968));
    CascadeMux I__2743 (
            .O(N__18977),
            .I(N__18965));
    InMux I__2742 (
            .O(N__18976),
            .I(N__18961));
    CascadeMux I__2741 (
            .O(N__18975),
            .I(N__18958));
    CascadeMux I__2740 (
            .O(N__18974),
            .I(N__18955));
    CascadeMux I__2739 (
            .O(N__18973),
            .I(N__18951));
    CascadeMux I__2738 (
            .O(N__18972),
            .I(N__18942));
    CascadeMux I__2737 (
            .O(N__18971),
            .I(N__18939));
    LocalMux I__2736 (
            .O(N__18968),
            .I(N__18936));
    InMux I__2735 (
            .O(N__18965),
            .I(N__18931));
    InMux I__2734 (
            .O(N__18964),
            .I(N__18931));
    LocalMux I__2733 (
            .O(N__18961),
            .I(N__18928));
    InMux I__2732 (
            .O(N__18958),
            .I(N__18925));
    InMux I__2731 (
            .O(N__18955),
            .I(N__18914));
    InMux I__2730 (
            .O(N__18954),
            .I(N__18914));
    InMux I__2729 (
            .O(N__18951),
            .I(N__18914));
    InMux I__2728 (
            .O(N__18950),
            .I(N__18914));
    InMux I__2727 (
            .O(N__18949),
            .I(N__18914));
    InMux I__2726 (
            .O(N__18948),
            .I(N__18901));
    InMux I__2725 (
            .O(N__18947),
            .I(N__18901));
    InMux I__2724 (
            .O(N__18946),
            .I(N__18901));
    InMux I__2723 (
            .O(N__18945),
            .I(N__18901));
    InMux I__2722 (
            .O(N__18942),
            .I(N__18901));
    InMux I__2721 (
            .O(N__18939),
            .I(N__18901));
    Odrv12 I__2720 (
            .O(N__18936),
            .I(\QuadInstance3.count_enable ));
    LocalMux I__2719 (
            .O(N__18931),
            .I(\QuadInstance3.count_enable ));
    Odrv4 I__2718 (
            .O(N__18928),
            .I(\QuadInstance3.count_enable ));
    LocalMux I__2717 (
            .O(N__18925),
            .I(\QuadInstance3.count_enable ));
    LocalMux I__2716 (
            .O(N__18914),
            .I(\QuadInstance3.count_enable ));
    LocalMux I__2715 (
            .O(N__18901),
            .I(\QuadInstance3.count_enable ));
    InMux I__2714 (
            .O(N__18888),
            .I(N__18885));
    LocalMux I__2713 (
            .O(N__18885),
            .I(N__18882));
    Odrv4 I__2712 (
            .O(N__18882),
            .I(\QuadInstance3.un1_Quad_axb_15 ));
    InMux I__2711 (
            .O(N__18879),
            .I(N__18876));
    LocalMux I__2710 (
            .O(N__18876),
            .I(N__18873));
    Span4Mux_v I__2709 (
            .O(N__18873),
            .I(N__18870));
    Span4Mux_v I__2708 (
            .O(N__18870),
            .I(N__18867));
    Odrv4 I__2707 (
            .O(N__18867),
            .I(\QuadInstance3.delayedCh_BZ0Z_0 ));
    InMux I__2706 (
            .O(N__18864),
            .I(N__18860));
    InMux I__2705 (
            .O(N__18863),
            .I(N__18857));
    LocalMux I__2704 (
            .O(N__18860),
            .I(\QuadInstance3.delayedCh_BZ0Z_1 ));
    LocalMux I__2703 (
            .O(N__18857),
            .I(\QuadInstance3.delayedCh_BZ0Z_1 ));
    InMux I__2702 (
            .O(N__18852),
            .I(\QuadInstance3.un1_Quad_cry_13 ));
    InMux I__2701 (
            .O(N__18849),
            .I(\QuadInstance3.un1_Quad_cry_14 ));
    CascadeMux I__2700 (
            .O(N__18846),
            .I(\QuadInstance3.count_enable_cascade_ ));
    CascadeMux I__2699 (
            .O(N__18843),
            .I(N__18840));
    InMux I__2698 (
            .O(N__18840),
            .I(N__18837));
    LocalMux I__2697 (
            .O(N__18837),
            .I(N__18834));
    Odrv4 I__2696 (
            .O(N__18834),
            .I(\QuadInstance3.Quad_RNI8OAL1Z0Z_1 ));
    CascadeMux I__2695 (
            .O(N__18831),
            .I(\QuadInstance3.un1_count_enable_i_a2_0_1_cascade_ ));
    CascadeMux I__2694 (
            .O(N__18828),
            .I(N__18825));
    InMux I__2693 (
            .O(N__18825),
            .I(N__18822));
    LocalMux I__2692 (
            .O(N__18822),
            .I(N__18819));
    Odrv4 I__2691 (
            .O(N__18819),
            .I(\QuadInstance3.Quad_RNI9PAL1Z0Z_2 ));
    CascadeMux I__2690 (
            .O(N__18816),
            .I(N__18813));
    InMux I__2689 (
            .O(N__18813),
            .I(N__18810));
    LocalMux I__2688 (
            .O(N__18810),
            .I(\QuadInstance3.Quad_RNIO10J1Z0Z_10 ));
    CascadeMux I__2687 (
            .O(N__18807),
            .I(N__18804));
    InMux I__2686 (
            .O(N__18804),
            .I(N__18801));
    LocalMux I__2685 (
            .O(N__18801),
            .I(\QuadInstance3.Quad_RNIFVAL1Z0Z_8 ));
    CascadeMux I__2684 (
            .O(N__18798),
            .I(N__18795));
    InMux I__2683 (
            .O(N__18795),
            .I(N__18792));
    LocalMux I__2682 (
            .O(N__18792),
            .I(\QuadInstance3.Quad_RNIG0BL1Z0Z_9 ));
    CascadeMux I__2681 (
            .O(N__18789),
            .I(N__18786));
    InMux I__2680 (
            .O(N__18786),
            .I(N__18783));
    LocalMux I__2679 (
            .O(N__18783),
            .I(N__18780));
    Odrv4 I__2678 (
            .O(N__18780),
            .I(\QuadInstance3.Quad_RNICSAL1Z0Z_5 ));
    InMux I__2677 (
            .O(N__18777),
            .I(\QuadInstance3.un1_Quad_cry_4 ));
    CascadeMux I__2676 (
            .O(N__18774),
            .I(N__18771));
    InMux I__2675 (
            .O(N__18771),
            .I(N__18768));
    LocalMux I__2674 (
            .O(N__18768),
            .I(N__18765));
    Odrv4 I__2673 (
            .O(N__18765),
            .I(\QuadInstance3.Quad_RNIDTAL1Z0Z_6 ));
    InMux I__2672 (
            .O(N__18762),
            .I(\QuadInstance3.un1_Quad_cry_5 ));
    InMux I__2671 (
            .O(N__18759),
            .I(\QuadInstance3.un1_Quad_cry_6 ));
    InMux I__2670 (
            .O(N__18756),
            .I(bfn_10_9_0_));
    InMux I__2669 (
            .O(N__18753),
            .I(\QuadInstance3.un1_Quad_cry_8 ));
    InMux I__2668 (
            .O(N__18750),
            .I(\QuadInstance3.un1_Quad_cry_9 ));
    CascadeMux I__2667 (
            .O(N__18747),
            .I(N__18744));
    InMux I__2666 (
            .O(N__18744),
            .I(N__18741));
    LocalMux I__2665 (
            .O(N__18741),
            .I(\QuadInstance3.Quad_RNIP20J1Z0Z_11 ));
    InMux I__2664 (
            .O(N__18738),
            .I(\QuadInstance3.un1_Quad_cry_10 ));
    CascadeMux I__2663 (
            .O(N__18735),
            .I(N__18732));
    InMux I__2662 (
            .O(N__18732),
            .I(N__18729));
    LocalMux I__2661 (
            .O(N__18729),
            .I(\QuadInstance3.Quad_RNIQ30J1Z0Z_12 ));
    InMux I__2660 (
            .O(N__18726),
            .I(\QuadInstance3.un1_Quad_cry_11 ));
    CascadeMux I__2659 (
            .O(N__18723),
            .I(N__18720));
    InMux I__2658 (
            .O(N__18720),
            .I(N__18717));
    LocalMux I__2657 (
            .O(N__18717),
            .I(\QuadInstance3.Quad_RNIR40J1Z0Z_13 ));
    InMux I__2656 (
            .O(N__18714),
            .I(\QuadInstance3.un1_Quad_cry_12 ));
    InMux I__2655 (
            .O(N__18711),
            .I(N__18708));
    LocalMux I__2654 (
            .O(N__18708),
            .I(\QuadInstance5.Quad_RNIBDQ82Z0Z_13 ));
    InMux I__2653 (
            .O(N__18705),
            .I(N__18702));
    LocalMux I__2652 (
            .O(N__18702),
            .I(\QuadInstance5.Quad_RNO_0_5_13 ));
    InMux I__2651 (
            .O(N__18699),
            .I(\QuadInstance5.un1_Quad_cry_12 ));
    InMux I__2650 (
            .O(N__18696),
            .I(N__18693));
    LocalMux I__2649 (
            .O(N__18693),
            .I(\QuadInstance5.Quad_RNICEQ82Z0Z_14 ));
    InMux I__2648 (
            .O(N__18690),
            .I(N__18687));
    LocalMux I__2647 (
            .O(N__18687),
            .I(\QuadInstance5.Quad_RNO_0_5_14 ));
    InMux I__2646 (
            .O(N__18684),
            .I(\QuadInstance5.un1_Quad_cry_13 ));
    InMux I__2645 (
            .O(N__18681),
            .I(N__18678));
    LocalMux I__2644 (
            .O(N__18678),
            .I(\QuadInstance5.un1_Quad_axb_15 ));
    InMux I__2643 (
            .O(N__18675),
            .I(\QuadInstance5.un1_Quad_cry_14 ));
    InMux I__2642 (
            .O(N__18672),
            .I(\QuadInstance3.un1_Quad_cry_0 ));
    InMux I__2641 (
            .O(N__18669),
            .I(\QuadInstance3.un1_Quad_cry_1 ));
    CascadeMux I__2640 (
            .O(N__18666),
            .I(N__18663));
    InMux I__2639 (
            .O(N__18663),
            .I(N__18660));
    LocalMux I__2638 (
            .O(N__18660),
            .I(N__18657));
    Odrv4 I__2637 (
            .O(N__18657),
            .I(\QuadInstance3.Quad_RNIAQAL1Z0Z_3 ));
    InMux I__2636 (
            .O(N__18654),
            .I(\QuadInstance3.un1_Quad_cry_2 ));
    InMux I__2635 (
            .O(N__18651),
            .I(\QuadInstance3.un1_Quad_cry_3 ));
    CascadeMux I__2634 (
            .O(N__18648),
            .I(N__18645));
    InMux I__2633 (
            .O(N__18645),
            .I(N__18642));
    LocalMux I__2632 (
            .O(N__18642),
            .I(\QuadInstance5.Quad_RNIR1LI2Z0Z_4 ));
    InMux I__2631 (
            .O(N__18639),
            .I(\QuadInstance5.un1_Quad_cry_3 ));
    CascadeMux I__2630 (
            .O(N__18636),
            .I(N__18633));
    InMux I__2629 (
            .O(N__18633),
            .I(N__18630));
    LocalMux I__2628 (
            .O(N__18630),
            .I(\QuadInstance5.Quad_RNIS2LI2Z0Z_5 ));
    InMux I__2627 (
            .O(N__18627),
            .I(\QuadInstance5.un1_Quad_cry_4 ));
    CascadeMux I__2626 (
            .O(N__18624),
            .I(N__18621));
    InMux I__2625 (
            .O(N__18621),
            .I(N__18618));
    LocalMux I__2624 (
            .O(N__18618),
            .I(\QuadInstance5.Quad_RNIT3LI2Z0Z_6 ));
    InMux I__2623 (
            .O(N__18615),
            .I(\QuadInstance5.un1_Quad_cry_5 ));
    InMux I__2622 (
            .O(N__18612),
            .I(N__18609));
    LocalMux I__2621 (
            .O(N__18609),
            .I(\QuadInstance5.Quad_RNIU4LI2Z0Z_7 ));
    InMux I__2620 (
            .O(N__18606),
            .I(\QuadInstance5.un1_Quad_cry_6 ));
    CascadeMux I__2619 (
            .O(N__18603),
            .I(N__18600));
    InMux I__2618 (
            .O(N__18600),
            .I(N__18597));
    LocalMux I__2617 (
            .O(N__18597),
            .I(\QuadInstance5.Quad_RNIV5LI2Z0Z_8 ));
    InMux I__2616 (
            .O(N__18594),
            .I(bfn_10_7_0_));
    CascadeMux I__2615 (
            .O(N__18591),
            .I(N__18588));
    InMux I__2614 (
            .O(N__18588),
            .I(N__18585));
    LocalMux I__2613 (
            .O(N__18585),
            .I(N__18582));
    Odrv4 I__2612 (
            .O(N__18582),
            .I(\QuadInstance5.Quad_RNI07LI2Z0Z_9 ));
    InMux I__2611 (
            .O(N__18579),
            .I(\QuadInstance5.un1_Quad_cry_8 ));
    CascadeMux I__2610 (
            .O(N__18576),
            .I(N__18573));
    InMux I__2609 (
            .O(N__18573),
            .I(N__18570));
    LocalMux I__2608 (
            .O(N__18570),
            .I(\QuadInstance5.Quad_RNI8AQ82Z0Z_10 ));
    InMux I__2607 (
            .O(N__18567),
            .I(\QuadInstance5.un1_Quad_cry_9 ));
    CascadeMux I__2606 (
            .O(N__18564),
            .I(N__18561));
    InMux I__2605 (
            .O(N__18561),
            .I(N__18558));
    LocalMux I__2604 (
            .O(N__18558),
            .I(\QuadInstance5.Quad_RNI9BQ82Z0Z_11 ));
    InMux I__2603 (
            .O(N__18555),
            .I(\QuadInstance5.un1_Quad_cry_10 ));
    CascadeMux I__2602 (
            .O(N__18552),
            .I(N__18549));
    InMux I__2601 (
            .O(N__18549),
            .I(N__18546));
    LocalMux I__2600 (
            .O(N__18546),
            .I(\QuadInstance5.Quad_RNIACQ82Z0Z_12 ));
    InMux I__2599 (
            .O(N__18543),
            .I(N__18540));
    LocalMux I__2598 (
            .O(N__18540),
            .I(\QuadInstance5.Quad_RNO_0_5_12 ));
    InMux I__2597 (
            .O(N__18537),
            .I(\QuadInstance5.un1_Quad_cry_11 ));
    InMux I__2596 (
            .O(N__18534),
            .I(N__18531));
    LocalMux I__2595 (
            .O(N__18531),
            .I(N__18526));
    InMux I__2594 (
            .O(N__18530),
            .I(N__18523));
    InMux I__2593 (
            .O(N__18529),
            .I(N__18520));
    Span4Mux_v I__2592 (
            .O(N__18526),
            .I(N__18508));
    LocalMux I__2591 (
            .O(N__18523),
            .I(N__18508));
    LocalMux I__2590 (
            .O(N__18520),
            .I(N__18508));
    CascadeMux I__2589 (
            .O(N__18519),
            .I(N__18500));
    CascadeMux I__2588 (
            .O(N__18518),
            .I(N__18496));
    CascadeMux I__2587 (
            .O(N__18517),
            .I(N__18493));
    CascadeMux I__2586 (
            .O(N__18516),
            .I(N__18488));
    InMux I__2585 (
            .O(N__18515),
            .I(N__18485));
    Span4Mux_h I__2584 (
            .O(N__18508),
            .I(N__18482));
    InMux I__2583 (
            .O(N__18507),
            .I(N__18473));
    InMux I__2582 (
            .O(N__18506),
            .I(N__18473));
    InMux I__2581 (
            .O(N__18505),
            .I(N__18473));
    InMux I__2580 (
            .O(N__18504),
            .I(N__18473));
    InMux I__2579 (
            .O(N__18503),
            .I(N__18456));
    InMux I__2578 (
            .O(N__18500),
            .I(N__18456));
    InMux I__2577 (
            .O(N__18499),
            .I(N__18456));
    InMux I__2576 (
            .O(N__18496),
            .I(N__18456));
    InMux I__2575 (
            .O(N__18493),
            .I(N__18456));
    InMux I__2574 (
            .O(N__18492),
            .I(N__18456));
    InMux I__2573 (
            .O(N__18491),
            .I(N__18456));
    InMux I__2572 (
            .O(N__18488),
            .I(N__18456));
    LocalMux I__2571 (
            .O(N__18485),
            .I(\QuadInstance2.count_enable ));
    Odrv4 I__2570 (
            .O(N__18482),
            .I(\QuadInstance2.count_enable ));
    LocalMux I__2569 (
            .O(N__18473),
            .I(\QuadInstance2.count_enable ));
    LocalMux I__2568 (
            .O(N__18456),
            .I(\QuadInstance2.count_enable ));
    InMux I__2567 (
            .O(N__18447),
            .I(N__18443));
    InMux I__2566 (
            .O(N__18446),
            .I(N__18440));
    LocalMux I__2565 (
            .O(N__18443),
            .I(\QuadInstance5.delayedCh_BZ0Z_1 ));
    LocalMux I__2564 (
            .O(N__18440),
            .I(\QuadInstance5.delayedCh_BZ0Z_1 ));
    InMux I__2563 (
            .O(N__18435),
            .I(N__18430));
    InMux I__2562 (
            .O(N__18434),
            .I(N__18427));
    InMux I__2561 (
            .O(N__18433),
            .I(N__18424));
    LocalMux I__2560 (
            .O(N__18430),
            .I(\QuadInstance5.delayedCh_AZ0Z_1 ));
    LocalMux I__2559 (
            .O(N__18427),
            .I(\QuadInstance5.delayedCh_AZ0Z_1 ));
    LocalMux I__2558 (
            .O(N__18424),
            .I(\QuadInstance5.delayedCh_AZ0Z_1 ));
    CascadeMux I__2557 (
            .O(N__18417),
            .I(N__18414));
    InMux I__2556 (
            .O(N__18414),
            .I(N__18411));
    LocalMux I__2555 (
            .O(N__18411),
            .I(\QuadInstance5.delayedCh_AZ0Z_2 ));
    InMux I__2554 (
            .O(N__18408),
            .I(N__18404));
    InMux I__2553 (
            .O(N__18407),
            .I(N__18401));
    LocalMux I__2552 (
            .O(N__18404),
            .I(\QuadInstance5.delayedCh_BZ0Z_2 ));
    LocalMux I__2551 (
            .O(N__18401),
            .I(\QuadInstance5.delayedCh_BZ0Z_2 ));
    CascadeMux I__2550 (
            .O(N__18396),
            .I(\QuadInstance5.count_enable_cascade_ ));
    CascadeMux I__2549 (
            .O(N__18393),
            .I(N__18389));
    CascadeMux I__2548 (
            .O(N__18392),
            .I(N__18384));
    InMux I__2547 (
            .O(N__18389),
            .I(N__18370));
    InMux I__2546 (
            .O(N__18388),
            .I(N__18370));
    InMux I__2545 (
            .O(N__18387),
            .I(N__18370));
    InMux I__2544 (
            .O(N__18384),
            .I(N__18370));
    CascadeMux I__2543 (
            .O(N__18383),
            .I(N__18365));
    CascadeMux I__2542 (
            .O(N__18382),
            .I(N__18361));
    CascadeMux I__2541 (
            .O(N__18381),
            .I(N__18355));
    CascadeMux I__2540 (
            .O(N__18380),
            .I(N__18352));
    CascadeMux I__2539 (
            .O(N__18379),
            .I(N__18348));
    LocalMux I__2538 (
            .O(N__18370),
            .I(N__18345));
    InMux I__2537 (
            .O(N__18369),
            .I(N__18342));
    InMux I__2536 (
            .O(N__18368),
            .I(N__18331));
    InMux I__2535 (
            .O(N__18365),
            .I(N__18331));
    InMux I__2534 (
            .O(N__18364),
            .I(N__18331));
    InMux I__2533 (
            .O(N__18361),
            .I(N__18331));
    InMux I__2532 (
            .O(N__18360),
            .I(N__18331));
    InMux I__2531 (
            .O(N__18359),
            .I(N__18318));
    InMux I__2530 (
            .O(N__18358),
            .I(N__18318));
    InMux I__2529 (
            .O(N__18355),
            .I(N__18318));
    InMux I__2528 (
            .O(N__18352),
            .I(N__18318));
    InMux I__2527 (
            .O(N__18351),
            .I(N__18318));
    InMux I__2526 (
            .O(N__18348),
            .I(N__18318));
    Odrv4 I__2525 (
            .O(N__18345),
            .I(\QuadInstance5.count_enable ));
    LocalMux I__2524 (
            .O(N__18342),
            .I(\QuadInstance5.count_enable ));
    LocalMux I__2523 (
            .O(N__18331),
            .I(\QuadInstance5.count_enable ));
    LocalMux I__2522 (
            .O(N__18318),
            .I(\QuadInstance5.count_enable ));
    CascadeMux I__2521 (
            .O(N__18309),
            .I(N__18306));
    InMux I__2520 (
            .O(N__18306),
            .I(N__18303));
    LocalMux I__2519 (
            .O(N__18303),
            .I(\QuadInstance5.Quad_RNIOUKI2Z0Z_1 ));
    InMux I__2518 (
            .O(N__18300),
            .I(N__18297));
    LocalMux I__2517 (
            .O(N__18297),
            .I(\QuadInstance5.Quad_RNO_0_4_1 ));
    InMux I__2516 (
            .O(N__18294),
            .I(\QuadInstance5.un1_Quad_cry_0 ));
    CascadeMux I__2515 (
            .O(N__18291),
            .I(N__18288));
    InMux I__2514 (
            .O(N__18288),
            .I(N__18285));
    LocalMux I__2513 (
            .O(N__18285),
            .I(\QuadInstance5.Quad_RNIPVKI2Z0Z_2 ));
    InMux I__2512 (
            .O(N__18282),
            .I(\QuadInstance5.un1_Quad_cry_1 ));
    CascadeMux I__2511 (
            .O(N__18279),
            .I(N__18276));
    InMux I__2510 (
            .O(N__18276),
            .I(N__18273));
    LocalMux I__2509 (
            .O(N__18273),
            .I(\QuadInstance5.Quad_RNIQ0LI2Z0Z_3 ));
    InMux I__2508 (
            .O(N__18270),
            .I(\QuadInstance5.un1_Quad_cry_2 ));
    InMux I__2507 (
            .O(N__18267),
            .I(N__18264));
    LocalMux I__2506 (
            .O(N__18264),
            .I(\PWMInstance0.PWMPulseWidthCountZ0Z_1 ));
    InMux I__2505 (
            .O(N__18261),
            .I(N__18258));
    LocalMux I__2504 (
            .O(N__18258),
            .I(N__18255));
    Span4Mux_h I__2503 (
            .O(N__18255),
            .I(N__18252));
    Odrv4 I__2502 (
            .O(N__18252),
            .I(\PWMInstance0.PWMPulseWidthCountZ0Z_7 ));
    CEMux I__2501 (
            .O(N__18249),
            .I(N__18245));
    CEMux I__2500 (
            .O(N__18248),
            .I(N__18242));
    LocalMux I__2499 (
            .O(N__18245),
            .I(N__18239));
    LocalMux I__2498 (
            .O(N__18242),
            .I(N__18236));
    Span4Mux_v I__2497 (
            .O(N__18239),
            .I(N__18228));
    Span4Mux_v I__2496 (
            .O(N__18236),
            .I(N__18228));
    CEMux I__2495 (
            .O(N__18235),
            .I(N__18225));
    CEMux I__2494 (
            .O(N__18234),
            .I(N__18222));
    CEMux I__2493 (
            .O(N__18233),
            .I(N__18219));
    Odrv4 I__2492 (
            .O(N__18228),
            .I(\PWMInstance0.pwmWrite_0_0 ));
    LocalMux I__2491 (
            .O(N__18225),
            .I(\PWMInstance0.pwmWrite_0_0 ));
    LocalMux I__2490 (
            .O(N__18222),
            .I(\PWMInstance0.pwmWrite_0_0 ));
    LocalMux I__2489 (
            .O(N__18219),
            .I(\PWMInstance0.pwmWrite_0_0 ));
    InMux I__2488 (
            .O(N__18210),
            .I(N__18207));
    LocalMux I__2487 (
            .O(N__18207),
            .I(N__18204));
    Odrv4 I__2486 (
            .O(N__18204),
            .I(\PWMInstance5.PWMPulseWidthCountZ0Z_13 ));
    InMux I__2485 (
            .O(N__18201),
            .I(N__18198));
    LocalMux I__2484 (
            .O(N__18198),
            .I(N__18195));
    Span12Mux_h I__2483 (
            .O(N__18195),
            .I(N__18192));
    Odrv12 I__2482 (
            .O(N__18192),
            .I(ch5_B_c));
    InMux I__2481 (
            .O(N__18189),
            .I(N__18186));
    LocalMux I__2480 (
            .O(N__18186),
            .I(N__18183));
    Odrv4 I__2479 (
            .O(N__18183),
            .I(\QuadInstance5.delayedCh_BZ0Z_0 ));
    InMux I__2478 (
            .O(N__18180),
            .I(\PWMInstance5.un1_periodCounter_2_cry_11 ));
    CascadeMux I__2477 (
            .O(N__18177),
            .I(N__18174));
    InMux I__2476 (
            .O(N__18174),
            .I(N__18169));
    InMux I__2475 (
            .O(N__18173),
            .I(N__18166));
    InMux I__2474 (
            .O(N__18172),
            .I(N__18163));
    LocalMux I__2473 (
            .O(N__18169),
            .I(N__18158));
    LocalMux I__2472 (
            .O(N__18166),
            .I(N__18158));
    LocalMux I__2471 (
            .O(N__18163),
            .I(\PWMInstance5.periodCounterZ0Z_13 ));
    Odrv4 I__2470 (
            .O(N__18158),
            .I(\PWMInstance5.periodCounterZ0Z_13 ));
    InMux I__2469 (
            .O(N__18153),
            .I(\PWMInstance5.un1_periodCounter_2_cry_12 ));
    InMux I__2468 (
            .O(N__18150),
            .I(\PWMInstance5.un1_periodCounter_2_cry_13 ));
    InMux I__2467 (
            .O(N__18147),
            .I(\PWMInstance5.un1_periodCounter_2_cry_14 ));
    InMux I__2466 (
            .O(N__18144),
            .I(bfn_9_14_0_));
    InMux I__2465 (
            .O(N__18141),
            .I(N__18137));
    InMux I__2464 (
            .O(N__18140),
            .I(N__18134));
    LocalMux I__2463 (
            .O(N__18137),
            .I(N__18130));
    LocalMux I__2462 (
            .O(N__18134),
            .I(N__18127));
    InMux I__2461 (
            .O(N__18133),
            .I(N__18124));
    Span4Mux_h I__2460 (
            .O(N__18130),
            .I(N__18121));
    Span4Mux_h I__2459 (
            .O(N__18127),
            .I(N__18118));
    LocalMux I__2458 (
            .O(N__18124),
            .I(\PWMInstance0.periodCounterZ0Z_8 ));
    Odrv4 I__2457 (
            .O(N__18121),
            .I(\PWMInstance0.periodCounterZ0Z_8 ));
    Odrv4 I__2456 (
            .O(N__18118),
            .I(\PWMInstance0.periodCounterZ0Z_8 ));
    CascadeMux I__2455 (
            .O(N__18111),
            .I(N__18107));
    InMux I__2454 (
            .O(N__18110),
            .I(N__18104));
    InMux I__2453 (
            .O(N__18107),
            .I(N__18101));
    LocalMux I__2452 (
            .O(N__18104),
            .I(N__18097));
    LocalMux I__2451 (
            .O(N__18101),
            .I(N__18094));
    InMux I__2450 (
            .O(N__18100),
            .I(N__18091));
    Span4Mux_h I__2449 (
            .O(N__18097),
            .I(N__18088));
    Span4Mux_h I__2448 (
            .O(N__18094),
            .I(N__18085));
    LocalMux I__2447 (
            .O(N__18091),
            .I(\PWMInstance0.periodCounterZ0Z_6 ));
    Odrv4 I__2446 (
            .O(N__18088),
            .I(\PWMInstance0.periodCounterZ0Z_6 ));
    Odrv4 I__2445 (
            .O(N__18085),
            .I(\PWMInstance0.periodCounterZ0Z_6 ));
    CascadeMux I__2444 (
            .O(N__18078),
            .I(N__18074));
    CascadeMux I__2443 (
            .O(N__18077),
            .I(N__18071));
    InMux I__2442 (
            .O(N__18074),
            .I(N__18068));
    InMux I__2441 (
            .O(N__18071),
            .I(N__18064));
    LocalMux I__2440 (
            .O(N__18068),
            .I(N__18061));
    InMux I__2439 (
            .O(N__18067),
            .I(N__18058));
    LocalMux I__2438 (
            .O(N__18064),
            .I(N__18055));
    Span4Mux_h I__2437 (
            .O(N__18061),
            .I(N__18052));
    LocalMux I__2436 (
            .O(N__18058),
            .I(\PWMInstance0.periodCounterZ0Z_13 ));
    Odrv4 I__2435 (
            .O(N__18055),
            .I(\PWMInstance0.periodCounterZ0Z_13 ));
    Odrv4 I__2434 (
            .O(N__18052),
            .I(\PWMInstance0.periodCounterZ0Z_13 ));
    InMux I__2433 (
            .O(N__18045),
            .I(N__18042));
    LocalMux I__2432 (
            .O(N__18042),
            .I(N__18039));
    Odrv4 I__2431 (
            .O(N__18039),
            .I(\PWMInstance0.un1_periodCounter12_1_0_a2_0_9 ));
    InMux I__2430 (
            .O(N__18036),
            .I(N__18029));
    InMux I__2429 (
            .O(N__18035),
            .I(N__18029));
    InMux I__2428 (
            .O(N__18034),
            .I(N__18026));
    LocalMux I__2427 (
            .O(N__18029),
            .I(N__18023));
    LocalMux I__2426 (
            .O(N__18026),
            .I(N__18018));
    Span4Mux_v I__2425 (
            .O(N__18023),
            .I(N__18018));
    Odrv4 I__2424 (
            .O(N__18018),
            .I(\PWMInstance0.periodCounterZ0Z_0 ));
    CascadeMux I__2423 (
            .O(N__18015),
            .I(N__18012));
    InMux I__2422 (
            .O(N__18012),
            .I(N__18008));
    InMux I__2421 (
            .O(N__18011),
            .I(N__18004));
    LocalMux I__2420 (
            .O(N__18008),
            .I(N__18001));
    InMux I__2419 (
            .O(N__18007),
            .I(N__17998));
    LocalMux I__2418 (
            .O(N__18004),
            .I(N__17993));
    Span4Mux_v I__2417 (
            .O(N__18001),
            .I(N__17993));
    LocalMux I__2416 (
            .O(N__17998),
            .I(\PWMInstance0.periodCounterZ0Z_1 ));
    Odrv4 I__2415 (
            .O(N__17993),
            .I(\PWMInstance0.periodCounterZ0Z_1 ));
    InMux I__2414 (
            .O(N__17988),
            .I(N__17985));
    LocalMux I__2413 (
            .O(N__17985),
            .I(\PWMInstance0.un1_PWMPulseWidthCount_0_I_1_c_RNOZ0 ));
    InMux I__2412 (
            .O(N__17982),
            .I(N__17979));
    LocalMux I__2411 (
            .O(N__17979),
            .I(\PWMInstance0.PWMPulseWidthCountZ0Z_0 ));
    InMux I__2410 (
            .O(N__17976),
            .I(\PWMInstance5.un1_periodCounter_2_cry_2 ));
    InMux I__2409 (
            .O(N__17973),
            .I(\PWMInstance5.un1_periodCounter_2_cry_3 ));
    InMux I__2408 (
            .O(N__17970),
            .I(\PWMInstance5.un1_periodCounter_2_cry_4 ));
    CascadeMux I__2407 (
            .O(N__17967),
            .I(N__17963));
    InMux I__2406 (
            .O(N__17966),
            .I(N__17959));
    InMux I__2405 (
            .O(N__17963),
            .I(N__17954));
    InMux I__2404 (
            .O(N__17962),
            .I(N__17954));
    LocalMux I__2403 (
            .O(N__17959),
            .I(\PWMInstance5.periodCounterZ0Z_6 ));
    LocalMux I__2402 (
            .O(N__17954),
            .I(\PWMInstance5.periodCounterZ0Z_6 ));
    InMux I__2401 (
            .O(N__17949),
            .I(\PWMInstance5.un1_periodCounter_2_cry_5 ));
    InMux I__2400 (
            .O(N__17946),
            .I(\PWMInstance5.un1_periodCounter_2_cry_6 ));
    InMux I__2399 (
            .O(N__17943),
            .I(N__17938));
    InMux I__2398 (
            .O(N__17942),
            .I(N__17935));
    InMux I__2397 (
            .O(N__17941),
            .I(N__17932));
    LocalMux I__2396 (
            .O(N__17938),
            .I(N__17929));
    LocalMux I__2395 (
            .O(N__17935),
            .I(N__17926));
    LocalMux I__2394 (
            .O(N__17932),
            .I(\PWMInstance5.periodCounterZ0Z_8 ));
    Odrv4 I__2393 (
            .O(N__17929),
            .I(\PWMInstance5.periodCounterZ0Z_8 ));
    Odrv12 I__2392 (
            .O(N__17926),
            .I(\PWMInstance5.periodCounterZ0Z_8 ));
    InMux I__2391 (
            .O(N__17919),
            .I(bfn_9_13_0_));
    InMux I__2390 (
            .O(N__17916),
            .I(\PWMInstance5.un1_periodCounter_2_cry_8 ));
    InMux I__2389 (
            .O(N__17913),
            .I(\PWMInstance5.un1_periodCounter_2_cry_9 ));
    InMux I__2388 (
            .O(N__17910),
            .I(\PWMInstance5.un1_periodCounter_2_cry_10 ));
    InMux I__2387 (
            .O(N__17907),
            .I(N__17904));
    LocalMux I__2386 (
            .O(N__17904),
            .I(N__17901));
    Span4Mux_v I__2385 (
            .O(N__17901),
            .I(N__17898));
    Odrv4 I__2384 (
            .O(N__17898),
            .I(\PWMInstance5.un1_PWMPulseWidthCount_0_I_1_c_RNO_4 ));
    InMux I__2383 (
            .O(N__17895),
            .I(N__17892));
    LocalMux I__2382 (
            .O(N__17892),
            .I(\PWMInstance5.PWMPulseWidthCountZ0Z_0 ));
    InMux I__2381 (
            .O(N__17889),
            .I(N__17886));
    LocalMux I__2380 (
            .O(N__17886),
            .I(\PWMInstance5.PWMPulseWidthCountZ0Z_1 ));
    InMux I__2379 (
            .O(N__17883),
            .I(N__17880));
    LocalMux I__2378 (
            .O(N__17880),
            .I(N__17877));
    Sp12to4 I__2377 (
            .O(N__17877),
            .I(N__17874));
    Odrv12 I__2376 (
            .O(N__17874),
            .I(\PWMInstance5.un1_PWMPulseWidthCount_0_I_27_c_RNO_4 ));
    InMux I__2375 (
            .O(N__17871),
            .I(N__17868));
    LocalMux I__2374 (
            .O(N__17868),
            .I(\PWMInstance5.PWMPulseWidthCountZ0Z_6 ));
    CascadeMux I__2373 (
            .O(N__17865),
            .I(N__17862));
    InMux I__2372 (
            .O(N__17862),
            .I(N__17859));
    LocalMux I__2371 (
            .O(N__17859),
            .I(\PWMInstance5.PWMPulseWidthCountZ0Z_7 ));
    InMux I__2370 (
            .O(N__17856),
            .I(N__17851));
    InMux I__2369 (
            .O(N__17855),
            .I(N__17846));
    InMux I__2368 (
            .O(N__17854),
            .I(N__17846));
    LocalMux I__2367 (
            .O(N__17851),
            .I(\PWMInstance5.periodCounterZ0Z_0 ));
    LocalMux I__2366 (
            .O(N__17846),
            .I(\PWMInstance5.periodCounterZ0Z_0 ));
    InMux I__2365 (
            .O(N__17841),
            .I(\PWMInstance5.un1_periodCounter_2_cry_0 ));
    InMux I__2364 (
            .O(N__17838),
            .I(\PWMInstance5.un1_periodCounter_2_cry_1 ));
    InMux I__2363 (
            .O(N__17835),
            .I(N__17832));
    LocalMux I__2362 (
            .O(N__17832),
            .I(N__17829));
    Odrv12 I__2361 (
            .O(N__17829),
            .I(\QuadInstance7.un1_Quad_axb_15 ));
    InMux I__2360 (
            .O(N__17826),
            .I(\QuadInstance7.un1_Quad_cry_14 ));
    InMux I__2359 (
            .O(N__17823),
            .I(N__17817));
    InMux I__2358 (
            .O(N__17822),
            .I(N__17817));
    LocalMux I__2357 (
            .O(N__17817),
            .I(pwmWrite_fastZ0Z_1));
    InMux I__2356 (
            .O(N__17814),
            .I(N__17808));
    InMux I__2355 (
            .O(N__17813),
            .I(N__17808));
    LocalMux I__2354 (
            .O(N__17808),
            .I(N__17804));
    InMux I__2353 (
            .O(N__17807),
            .I(N__17801));
    Span4Mux_h I__2352 (
            .O(N__17804),
            .I(N__17798));
    LocalMux I__2351 (
            .O(N__17801),
            .I(N__17795));
    Span4Mux_h I__2350 (
            .O(N__17798),
            .I(N__17792));
    Span4Mux_h I__2349 (
            .O(N__17795),
            .I(N__17789));
    Odrv4 I__2348 (
            .O(N__17792),
            .I(pwmWriteZ0Z_7));
    Odrv4 I__2347 (
            .O(N__17789),
            .I(pwmWriteZ0Z_7));
    CascadeMux I__2346 (
            .O(N__17784),
            .I(N__17781));
    InMux I__2345 (
            .O(N__17781),
            .I(N__17778));
    LocalMux I__2344 (
            .O(N__17778),
            .I(\QuadInstance7.Quad_RNIEBVV2Z0Z_7 ));
    InMux I__2343 (
            .O(N__17775),
            .I(\QuadInstance7.un1_Quad_cry_6 ));
    CascadeMux I__2342 (
            .O(N__17772),
            .I(N__17769));
    InMux I__2341 (
            .O(N__17769),
            .I(N__17766));
    LocalMux I__2340 (
            .O(N__17766),
            .I(\QuadInstance7.Quad_RNIFCVV2Z0Z_8 ));
    InMux I__2339 (
            .O(N__17763),
            .I(bfn_9_9_0_));
    CascadeMux I__2338 (
            .O(N__17760),
            .I(N__17757));
    InMux I__2337 (
            .O(N__17757),
            .I(N__17754));
    LocalMux I__2336 (
            .O(N__17754),
            .I(\QuadInstance7.Quad_RNIGDVV2Z0Z_9 ));
    InMux I__2335 (
            .O(N__17751),
            .I(\QuadInstance7.un1_Quad_cry_8 ));
    CascadeMux I__2334 (
            .O(N__17748),
            .I(N__17745));
    InMux I__2333 (
            .O(N__17745),
            .I(N__17742));
    LocalMux I__2332 (
            .O(N__17742),
            .I(\QuadInstance7.Quad_RNIOIKU2Z0Z_10 ));
    InMux I__2331 (
            .O(N__17739),
            .I(\QuadInstance7.un1_Quad_cry_9 ));
    CascadeMux I__2330 (
            .O(N__17736),
            .I(N__17733));
    InMux I__2329 (
            .O(N__17733),
            .I(N__17730));
    LocalMux I__2328 (
            .O(N__17730),
            .I(\QuadInstance7.Quad_RNIPJKU2Z0Z_11 ));
    InMux I__2327 (
            .O(N__17727),
            .I(N__17724));
    LocalMux I__2326 (
            .O(N__17724),
            .I(N__17721));
    Odrv4 I__2325 (
            .O(N__17721),
            .I(\QuadInstance7.Quad_RNO_0_7_11 ));
    InMux I__2324 (
            .O(N__17718),
            .I(\QuadInstance7.un1_Quad_cry_10 ));
    CascadeMux I__2323 (
            .O(N__17715),
            .I(N__17712));
    InMux I__2322 (
            .O(N__17712),
            .I(N__17709));
    LocalMux I__2321 (
            .O(N__17709),
            .I(\QuadInstance7.Quad_RNIQKKU2Z0Z_12 ));
    InMux I__2320 (
            .O(N__17706),
            .I(N__17703));
    LocalMux I__2319 (
            .O(N__17703),
            .I(N__17700));
    Odrv4 I__2318 (
            .O(N__17700),
            .I(\QuadInstance7.Quad_RNO_0_7_12 ));
    InMux I__2317 (
            .O(N__17697),
            .I(\QuadInstance7.un1_Quad_cry_11 ));
    CascadeMux I__2316 (
            .O(N__17694),
            .I(N__17691));
    InMux I__2315 (
            .O(N__17691),
            .I(N__17688));
    LocalMux I__2314 (
            .O(N__17688),
            .I(\QuadInstance7.Quad_RNIRLKU2Z0Z_13 ));
    InMux I__2313 (
            .O(N__17685),
            .I(\QuadInstance7.un1_Quad_cry_12 ));
    InMux I__2312 (
            .O(N__17682),
            .I(N__17679));
    LocalMux I__2311 (
            .O(N__17679),
            .I(\QuadInstance7.Quad_RNISMKU2Z0Z_14 ));
    InMux I__2310 (
            .O(N__17676),
            .I(\QuadInstance7.un1_Quad_cry_13 ));
    CascadeMux I__2309 (
            .O(N__17673),
            .I(N__17670));
    InMux I__2308 (
            .O(N__17670),
            .I(N__17667));
    LocalMux I__2307 (
            .O(N__17667),
            .I(\QuadInstance7.Quad_RNI85VV2Z0Z_1 ));
    InMux I__2306 (
            .O(N__17664),
            .I(\QuadInstance7.un1_Quad_cry_0 ));
    CascadeMux I__2305 (
            .O(N__17661),
            .I(N__17658));
    InMux I__2304 (
            .O(N__17658),
            .I(N__17655));
    LocalMux I__2303 (
            .O(N__17655),
            .I(\QuadInstance7.Quad_RNI96VV2Z0Z_2 ));
    InMux I__2302 (
            .O(N__17652),
            .I(\QuadInstance7.un1_Quad_cry_1 ));
    CascadeMux I__2301 (
            .O(N__17649),
            .I(N__17646));
    InMux I__2300 (
            .O(N__17646),
            .I(N__17643));
    LocalMux I__2299 (
            .O(N__17643),
            .I(\QuadInstance7.Quad_RNIA7VV2Z0Z_3 ));
    InMux I__2298 (
            .O(N__17640),
            .I(\QuadInstance7.un1_Quad_cry_2 ));
    CascadeMux I__2297 (
            .O(N__17637),
            .I(N__17634));
    InMux I__2296 (
            .O(N__17634),
            .I(N__17631));
    LocalMux I__2295 (
            .O(N__17631),
            .I(\QuadInstance7.Quad_RNIB8VV2Z0Z_4 ));
    InMux I__2294 (
            .O(N__17628),
            .I(\QuadInstance7.un1_Quad_cry_3 ));
    CascadeMux I__2293 (
            .O(N__17625),
            .I(N__17622));
    InMux I__2292 (
            .O(N__17622),
            .I(N__17619));
    LocalMux I__2291 (
            .O(N__17619),
            .I(\QuadInstance7.Quad_RNIC9VV2Z0Z_5 ));
    InMux I__2290 (
            .O(N__17616),
            .I(\QuadInstance7.un1_Quad_cry_4 ));
    CascadeMux I__2289 (
            .O(N__17613),
            .I(N__17610));
    InMux I__2288 (
            .O(N__17610),
            .I(N__17607));
    LocalMux I__2287 (
            .O(N__17607),
            .I(\QuadInstance7.Quad_RNIDAVV2Z0Z_6 ));
    InMux I__2286 (
            .O(N__17604),
            .I(\QuadInstance7.un1_Quad_cry_5 ));
    CascadeMux I__2285 (
            .O(N__17601),
            .I(N__17598));
    InMux I__2284 (
            .O(N__17598),
            .I(N__17595));
    LocalMux I__2283 (
            .O(N__17595),
            .I(N__17585));
    CascadeMux I__2282 (
            .O(N__17594),
            .I(N__17581));
    CascadeMux I__2281 (
            .O(N__17593),
            .I(N__17578));
    CascadeMux I__2280 (
            .O(N__17592),
            .I(N__17573));
    CascadeMux I__2279 (
            .O(N__17591),
            .I(N__17569));
    CascadeMux I__2278 (
            .O(N__17590),
            .I(N__17565));
    CascadeMux I__2277 (
            .O(N__17589),
            .I(N__17562));
    InMux I__2276 (
            .O(N__17588),
            .I(N__17558));
    Span4Mux_h I__2275 (
            .O(N__17585),
            .I(N__17555));
    InMux I__2274 (
            .O(N__17584),
            .I(N__17546));
    InMux I__2273 (
            .O(N__17581),
            .I(N__17546));
    InMux I__2272 (
            .O(N__17578),
            .I(N__17546));
    InMux I__2271 (
            .O(N__17577),
            .I(N__17546));
    InMux I__2270 (
            .O(N__17576),
            .I(N__17529));
    InMux I__2269 (
            .O(N__17573),
            .I(N__17529));
    InMux I__2268 (
            .O(N__17572),
            .I(N__17529));
    InMux I__2267 (
            .O(N__17569),
            .I(N__17529));
    InMux I__2266 (
            .O(N__17568),
            .I(N__17529));
    InMux I__2265 (
            .O(N__17565),
            .I(N__17529));
    InMux I__2264 (
            .O(N__17562),
            .I(N__17529));
    InMux I__2263 (
            .O(N__17561),
            .I(N__17529));
    LocalMux I__2262 (
            .O(N__17558),
            .I(\QuadInstance2.un1_count_enable_i_a2_0_1 ));
    Odrv4 I__2261 (
            .O(N__17555),
            .I(\QuadInstance2.un1_count_enable_i_a2_0_1 ));
    LocalMux I__2260 (
            .O(N__17546),
            .I(\QuadInstance2.un1_count_enable_i_a2_0_1 ));
    LocalMux I__2259 (
            .O(N__17529),
            .I(\QuadInstance2.un1_count_enable_i_a2_0_1 ));
    CascadeMux I__2258 (
            .O(N__17520),
            .I(N__17517));
    InMux I__2257 (
            .O(N__17517),
            .I(N__17514));
    LocalMux I__2256 (
            .O(N__17514),
            .I(N__17511));
    Span4Mux_h I__2255 (
            .O(N__17511),
            .I(N__17508));
    Odrv4 I__2254 (
            .O(N__17508),
            .I(\QuadInstance2.Quad_RNIJ03G2Z0Z_13 ));
    InMux I__2253 (
            .O(N__17505),
            .I(N__17490));
    InMux I__2252 (
            .O(N__17504),
            .I(N__17490));
    InMux I__2251 (
            .O(N__17503),
            .I(N__17490));
    InMux I__2250 (
            .O(N__17502),
            .I(N__17490));
    CascadeMux I__2249 (
            .O(N__17501),
            .I(N__17487));
    CascadeMux I__2248 (
            .O(N__17500),
            .I(N__17483));
    CascadeMux I__2247 (
            .O(N__17499),
            .I(N__17479));
    LocalMux I__2246 (
            .O(N__17490),
            .I(N__17471));
    InMux I__2245 (
            .O(N__17487),
            .I(N__17466));
    InMux I__2244 (
            .O(N__17486),
            .I(N__17466));
    InMux I__2243 (
            .O(N__17483),
            .I(N__17457));
    InMux I__2242 (
            .O(N__17482),
            .I(N__17457));
    InMux I__2241 (
            .O(N__17479),
            .I(N__17457));
    InMux I__2240 (
            .O(N__17478),
            .I(N__17457));
    InMux I__2239 (
            .O(N__17477),
            .I(N__17448));
    InMux I__2238 (
            .O(N__17476),
            .I(N__17448));
    InMux I__2237 (
            .O(N__17475),
            .I(N__17448));
    InMux I__2236 (
            .O(N__17474),
            .I(N__17448));
    Odrv4 I__2235 (
            .O(N__17471),
            .I(\QuadInstance5.un1_count_enable_i_a2_0_1 ));
    LocalMux I__2234 (
            .O(N__17466),
            .I(\QuadInstance5.un1_count_enable_i_a2_0_1 ));
    LocalMux I__2233 (
            .O(N__17457),
            .I(\QuadInstance5.un1_count_enable_i_a2_0_1 ));
    LocalMux I__2232 (
            .O(N__17448),
            .I(\QuadInstance5.un1_count_enable_i_a2_0_1 ));
    CascadeMux I__2231 (
            .O(N__17439),
            .I(\QuadInstance5.un1_count_enable_i_a2_0_1_cascade_ ));
    InMux I__2230 (
            .O(N__17436),
            .I(N__17433));
    LocalMux I__2229 (
            .O(N__17433),
            .I(N__17430));
    Span4Mux_h I__2228 (
            .O(N__17430),
            .I(N__17427));
    Span4Mux_h I__2227 (
            .O(N__17427),
            .I(N__17424));
    Span4Mux_h I__2226 (
            .O(N__17424),
            .I(N__17421));
    Odrv4 I__2225 (
            .O(N__17421),
            .I(ch7_B_c));
    InMux I__2224 (
            .O(N__17418),
            .I(N__17415));
    LocalMux I__2223 (
            .O(N__17415),
            .I(N__17412));
    Odrv12 I__2222 (
            .O(N__17412),
            .I(\QuadInstance7.delayedCh_BZ0Z_0 ));
    IoInMux I__2221 (
            .O(N__17409),
            .I(N__17406));
    LocalMux I__2220 (
            .O(N__17406),
            .I(PWM0_obufLegalizeSB_DFFNet));
    IoInMux I__2219 (
            .O(N__17403),
            .I(N__17400));
    LocalMux I__2218 (
            .O(N__17400),
            .I(PWM1_obufLegalizeSB_DFFNet));
    IoInMux I__2217 (
            .O(N__17397),
            .I(N__17394));
    LocalMux I__2216 (
            .O(N__17394),
            .I(PWM6_obufLegalizeSB_DFFNet));
    IoInMux I__2215 (
            .O(N__17391),
            .I(N__17388));
    LocalMux I__2214 (
            .O(N__17388),
            .I(PWM7_obufLegalizeSB_DFFNet));
    InMux I__2213 (
            .O(N__17385),
            .I(N__17382));
    LocalMux I__2212 (
            .O(N__17382),
            .I(N__17379));
    Odrv4 I__2211 (
            .O(N__17379),
            .I(ch3_B_c));
    InMux I__2210 (
            .O(N__17376),
            .I(N__17373));
    LocalMux I__2209 (
            .O(N__17373),
            .I(N__17370));
    Span4Mux_v I__2208 (
            .O(N__17370),
            .I(N__17367));
    Odrv4 I__2207 (
            .O(N__17367),
            .I(\QuadInstance2.Quad_RNO_0_2_4 ));
    InMux I__2206 (
            .O(N__17364),
            .I(N__17361));
    LocalMux I__2205 (
            .O(N__17361),
            .I(N__17358));
    Span4Mux_h I__2204 (
            .O(N__17358),
            .I(N__17355));
    Odrv4 I__2203 (
            .O(N__17355),
            .I(ch5_A_c));
    InMux I__2202 (
            .O(N__17352),
            .I(N__17349));
    LocalMux I__2201 (
            .O(N__17349),
            .I(\QuadInstance5.delayedCh_AZ0Z_0 ));
    InMux I__2200 (
            .O(N__17346),
            .I(N__17343));
    LocalMux I__2199 (
            .O(N__17343),
            .I(\PWMInstance0.un1_PWMPulseWidthCount_0_I_9_c_RNOZ0 ));
    InMux I__2198 (
            .O(N__17340),
            .I(N__17337));
    LocalMux I__2197 (
            .O(N__17337),
            .I(\PWMInstance0.un1_PWMPulseWidthCount_0_I_15_c_RNOZ0 ));
    InMux I__2196 (
            .O(N__17334),
            .I(N__17331));
    LocalMux I__2195 (
            .O(N__17331),
            .I(N__17328));
    Odrv4 I__2194 (
            .O(N__17328),
            .I(\PWMInstance0.un1_PWMPulseWidthCount_0_I_27_c_RNOZ0 ));
    InMux I__2193 (
            .O(N__17325),
            .I(N__17322));
    LocalMux I__2192 (
            .O(N__17322),
            .I(N__17319));
    Odrv4 I__2191 (
            .O(N__17319),
            .I(\PWMInstance0.un1_PWMPulseWidthCount_0_I_45_c_RNOZ0 ));
    InMux I__2190 (
            .O(N__17316),
            .I(N__17313));
    LocalMux I__2189 (
            .O(N__17313),
            .I(\PWMInstance0.un1_PWMPulseWidthCount_0_I_33_c_RNOZ0 ));
    InMux I__2188 (
            .O(N__17310),
            .I(N__17307));
    LocalMux I__2187 (
            .O(N__17307),
            .I(\PWMInstance0.un1_PWMPulseWidthCount_0_I_39_c_RNOZ0 ));
    InMux I__2186 (
            .O(N__17304),
            .I(N__17301));
    LocalMux I__2185 (
            .O(N__17301),
            .I(\PWMInstance0.un1_PWMPulseWidthCount_0_I_21_c_RNOZ0 ));
    InMux I__2184 (
            .O(N__17298),
            .I(N__17295));
    LocalMux I__2183 (
            .O(N__17295),
            .I(\PWMInstance0.un1_periodCounter12_1_0_a2_0 ));
    CascadeMux I__2182 (
            .O(N__17292),
            .I(N__17285));
    InMux I__2181 (
            .O(N__17291),
            .I(N__17281));
    InMux I__2180 (
            .O(N__17290),
            .I(N__17278));
    InMux I__2179 (
            .O(N__17289),
            .I(N__17273));
    InMux I__2178 (
            .O(N__17288),
            .I(N__17273));
    InMux I__2177 (
            .O(N__17285),
            .I(N__17270));
    InMux I__2176 (
            .O(N__17284),
            .I(N__17267));
    LocalMux I__2175 (
            .O(N__17281),
            .I(N__17260));
    LocalMux I__2174 (
            .O(N__17278),
            .I(N__17260));
    LocalMux I__2173 (
            .O(N__17273),
            .I(N__17260));
    LocalMux I__2172 (
            .O(N__17270),
            .I(\PWMInstance0.out_0_sqmuxa ));
    LocalMux I__2171 (
            .O(N__17267),
            .I(\PWMInstance0.out_0_sqmuxa ));
    Odrv12 I__2170 (
            .O(N__17260),
            .I(\PWMInstance0.out_0_sqmuxa ));
    InMux I__2169 (
            .O(N__17253),
            .I(bfn_8_16_0_));
    IoInMux I__2168 (
            .O(N__17250),
            .I(N__17247));
    LocalMux I__2167 (
            .O(N__17247),
            .I(N__17244));
    Span4Mux_s2_v I__2166 (
            .O(N__17244),
            .I(N__17240));
    InMux I__2165 (
            .O(N__17243),
            .I(N__17237));
    Odrv4 I__2164 (
            .O(N__17240),
            .I(PWM0_c));
    LocalMux I__2163 (
            .O(N__17237),
            .I(PWM0_c));
    InMux I__2162 (
            .O(N__17232),
            .I(N__17229));
    LocalMux I__2161 (
            .O(N__17229),
            .I(N__17226));
    Span4Mux_h I__2160 (
            .O(N__17226),
            .I(N__17223));
    Odrv4 I__2159 (
            .O(N__17223),
            .I(\PWMInstance5.PWMPulseWidthCountZ0Z_12 ));
    InMux I__2158 (
            .O(N__17220),
            .I(N__17217));
    LocalMux I__2157 (
            .O(N__17217),
            .I(N__17214));
    Span12Mux_s4_v I__2156 (
            .O(N__17214),
            .I(N__17211));
    Odrv12 I__2155 (
            .O(N__17211),
            .I(\PWMInstance5.un1_PWMPulseWidthCount_0_I_39_c_RNO_4 ));
    InMux I__2154 (
            .O(N__17208),
            .I(N__17205));
    LocalMux I__2153 (
            .O(N__17205),
            .I(\PWMInstance0.PWMPulseWidthCountZ0Z_6 ));
    InMux I__2152 (
            .O(N__17202),
            .I(N__17199));
    LocalMux I__2151 (
            .O(N__17199),
            .I(N__17195));
    InMux I__2150 (
            .O(N__17198),
            .I(N__17191));
    Span4Mux_h I__2149 (
            .O(N__17195),
            .I(N__17188));
    InMux I__2148 (
            .O(N__17194),
            .I(N__17185));
    LocalMux I__2147 (
            .O(N__17191),
            .I(\PWMInstance0.periodCounterZ0Z_7 ));
    Odrv4 I__2146 (
            .O(N__17188),
            .I(\PWMInstance0.periodCounterZ0Z_7 ));
    LocalMux I__2145 (
            .O(N__17185),
            .I(\PWMInstance0.periodCounterZ0Z_7 ));
    CascadeMux I__2144 (
            .O(N__17178),
            .I(N__17175));
    InMux I__2143 (
            .O(N__17175),
            .I(N__17172));
    LocalMux I__2142 (
            .O(N__17172),
            .I(N__17167));
    InMux I__2141 (
            .O(N__17171),
            .I(N__17164));
    InMux I__2140 (
            .O(N__17170),
            .I(N__17161));
    Span4Mux_h I__2139 (
            .O(N__17167),
            .I(N__17156));
    LocalMux I__2138 (
            .O(N__17164),
            .I(N__17156));
    LocalMux I__2137 (
            .O(N__17161),
            .I(\PWMInstance0.periodCounterZ0Z_15 ));
    Odrv4 I__2136 (
            .O(N__17156),
            .I(\PWMInstance0.periodCounterZ0Z_15 ));
    InMux I__2135 (
            .O(N__17151),
            .I(N__17148));
    LocalMux I__2134 (
            .O(N__17148),
            .I(N__17143));
    InMux I__2133 (
            .O(N__17147),
            .I(N__17140));
    InMux I__2132 (
            .O(N__17146),
            .I(N__17137));
    Span4Mux_h I__2131 (
            .O(N__17143),
            .I(N__17134));
    LocalMux I__2130 (
            .O(N__17140),
            .I(N__17131));
    LocalMux I__2129 (
            .O(N__17137),
            .I(\PWMInstance0.periodCounterZ0Z_14 ));
    Odrv4 I__2128 (
            .O(N__17134),
            .I(\PWMInstance0.periodCounterZ0Z_14 ));
    Odrv12 I__2127 (
            .O(N__17131),
            .I(\PWMInstance0.periodCounterZ0Z_14 ));
    InMux I__2126 (
            .O(N__17124),
            .I(N__17121));
    LocalMux I__2125 (
            .O(N__17121),
            .I(\PWMInstance0.PWMPulseWidthCountZ0Z_14 ));
    InMux I__2124 (
            .O(N__17118),
            .I(N__17115));
    LocalMux I__2123 (
            .O(N__17115),
            .I(\PWMInstance0.PWMPulseWidthCountZ0Z_15 ));
    InMux I__2122 (
            .O(N__17112),
            .I(N__17107));
    InMux I__2121 (
            .O(N__17111),
            .I(N__17104));
    InMux I__2120 (
            .O(N__17110),
            .I(N__17101));
    LocalMux I__2119 (
            .O(N__17107),
            .I(N__17098));
    LocalMux I__2118 (
            .O(N__17104),
            .I(N__17095));
    LocalMux I__2117 (
            .O(N__17101),
            .I(\PWMInstance0.periodCounterZ0Z_10 ));
    Odrv4 I__2116 (
            .O(N__17098),
            .I(\PWMInstance0.periodCounterZ0Z_10 ));
    Odrv4 I__2115 (
            .O(N__17095),
            .I(\PWMInstance0.periodCounterZ0Z_10 ));
    CascadeMux I__2114 (
            .O(N__17088),
            .I(N__17084));
    CascadeMux I__2113 (
            .O(N__17087),
            .I(N__17081));
    InMux I__2112 (
            .O(N__17084),
            .I(N__17077));
    InMux I__2111 (
            .O(N__17081),
            .I(N__17074));
    InMux I__2110 (
            .O(N__17080),
            .I(N__17071));
    LocalMux I__2109 (
            .O(N__17077),
            .I(N__17068));
    LocalMux I__2108 (
            .O(N__17074),
            .I(N__17065));
    LocalMux I__2107 (
            .O(N__17071),
            .I(\PWMInstance0.periodCounterZ0Z_11 ));
    Odrv4 I__2106 (
            .O(N__17068),
            .I(\PWMInstance0.periodCounterZ0Z_11 ));
    Odrv4 I__2105 (
            .O(N__17065),
            .I(\PWMInstance0.periodCounterZ0Z_11 ));
    InMux I__2104 (
            .O(N__17058),
            .I(N__17055));
    LocalMux I__2103 (
            .O(N__17055),
            .I(N__17052));
    Span4Mux_h I__2102 (
            .O(N__17052),
            .I(N__17049));
    Odrv4 I__2101 (
            .O(N__17049),
            .I(\PWMInstance0.PWMPulseWidthCountZ0Z_10 ));
    InMux I__2100 (
            .O(N__17046),
            .I(N__17043));
    LocalMux I__2099 (
            .O(N__17043),
            .I(\PWMInstance0.PWMPulseWidthCountZ0Z_11 ));
    InMux I__2098 (
            .O(N__17040),
            .I(N__17037));
    LocalMux I__2097 (
            .O(N__17037),
            .I(\PWMInstance0.PWMPulseWidthCountZ0Z_13 ));
    InMux I__2096 (
            .O(N__17034),
            .I(N__17031));
    LocalMux I__2095 (
            .O(N__17031),
            .I(\PWMInstance0.PWMPulseWidthCountZ0Z_12 ));
    InMux I__2094 (
            .O(N__17028),
            .I(N__17023));
    InMux I__2093 (
            .O(N__17027),
            .I(N__17020));
    InMux I__2092 (
            .O(N__17026),
            .I(N__17017));
    LocalMux I__2091 (
            .O(N__17023),
            .I(N__17014));
    LocalMux I__2090 (
            .O(N__17020),
            .I(N__17011));
    LocalMux I__2089 (
            .O(N__17017),
            .I(\PWMInstance0.periodCounterZ0Z_12 ));
    Odrv4 I__2088 (
            .O(N__17014),
            .I(\PWMInstance0.periodCounterZ0Z_12 ));
    Odrv4 I__2087 (
            .O(N__17011),
            .I(\PWMInstance0.periodCounterZ0Z_12 ));
    InMux I__2086 (
            .O(N__17004),
            .I(N__16996));
    InMux I__2085 (
            .O(N__17003),
            .I(N__16991));
    InMux I__2084 (
            .O(N__17002),
            .I(N__16991));
    InMux I__2083 (
            .O(N__17001),
            .I(N__16988));
    InMux I__2082 (
            .O(N__17000),
            .I(N__16985));
    CascadeMux I__2081 (
            .O(N__16999),
            .I(N__16982));
    LocalMux I__2080 (
            .O(N__16996),
            .I(N__16973));
    LocalMux I__2079 (
            .O(N__16991),
            .I(N__16973));
    LocalMux I__2078 (
            .O(N__16988),
            .I(N__16973));
    LocalMux I__2077 (
            .O(N__16985),
            .I(N__16973));
    InMux I__2076 (
            .O(N__16982),
            .I(N__16970));
    Span12Mux_s5_v I__2075 (
            .O(N__16973),
            .I(N__16967));
    LocalMux I__2074 (
            .O(N__16970),
            .I(\PWMInstance1.out_0_sqmuxa ));
    Odrv12 I__2073 (
            .O(N__16967),
            .I(\PWMInstance1.out_0_sqmuxa ));
    InMux I__2072 (
            .O(N__16962),
            .I(N__16959));
    LocalMux I__2071 (
            .O(N__16959),
            .I(N__16956));
    Odrv12 I__2070 (
            .O(N__16956),
            .I(\PWMInstance5.un1_PWMPulseWidthCount_0_I_9_c_RNO_4 ));
    InMux I__2069 (
            .O(N__16953),
            .I(N__16950));
    LocalMux I__2068 (
            .O(N__16950),
            .I(\PWMInstance5.PWMPulseWidthCountZ0Z_2 ));
    InMux I__2067 (
            .O(N__16947),
            .I(N__16944));
    LocalMux I__2066 (
            .O(N__16944),
            .I(\PWMInstance5.PWMPulseWidthCountZ0Z_3 ));
    InMux I__2065 (
            .O(N__16941),
            .I(N__16938));
    LocalMux I__2064 (
            .O(N__16938),
            .I(N__16935));
    Odrv4 I__2063 (
            .O(N__16935),
            .I(\PWMInstance5.PWMPulseWidthCountZ0Z_14 ));
    InMux I__2062 (
            .O(N__16932),
            .I(N__16929));
    LocalMux I__2061 (
            .O(N__16929),
            .I(N__16926));
    Span12Mux_s3_v I__2060 (
            .O(N__16926),
            .I(N__16923));
    Odrv12 I__2059 (
            .O(N__16923),
            .I(\PWMInstance5.un1_PWMPulseWidthCount_0_I_21_c_RNO_4 ));
    InMux I__2058 (
            .O(N__16920),
            .I(N__16917));
    LocalMux I__2057 (
            .O(N__16917),
            .I(\PWMInstance5.PWMPulseWidthCountZ0Z_15 ));
    InMux I__2056 (
            .O(N__16914),
            .I(N__16911));
    LocalMux I__2055 (
            .O(N__16911),
            .I(\PWMInstance0.PWMPulseWidthCountZ0Z_9 ));
    CascadeMux I__2054 (
            .O(N__16908),
            .I(N__16905));
    InMux I__2053 (
            .O(N__16905),
            .I(N__16901));
    InMux I__2052 (
            .O(N__16904),
            .I(N__16897));
    LocalMux I__2051 (
            .O(N__16901),
            .I(N__16894));
    InMux I__2050 (
            .O(N__16900),
            .I(N__16891));
    LocalMux I__2049 (
            .O(N__16897),
            .I(N__16886));
    Span4Mux_h I__2048 (
            .O(N__16894),
            .I(N__16886));
    LocalMux I__2047 (
            .O(N__16891),
            .I(\PWMInstance0.periodCounterZ0Z_9 ));
    Odrv4 I__2046 (
            .O(N__16886),
            .I(\PWMInstance0.periodCounterZ0Z_9 ));
    InMux I__2045 (
            .O(N__16881),
            .I(N__16878));
    LocalMux I__2044 (
            .O(N__16878),
            .I(\PWMInstance0.PWMPulseWidthCountZ0Z_8 ));
    InMux I__2043 (
            .O(N__16875),
            .I(N__16869));
    InMux I__2042 (
            .O(N__16874),
            .I(N__16869));
    LocalMux I__2041 (
            .O(N__16869),
            .I(N__16866));
    Span4Mux_h I__2040 (
            .O(N__16866),
            .I(N__16862));
    InMux I__2039 (
            .O(N__16865),
            .I(N__16859));
    Odrv4 I__2038 (
            .O(N__16862),
            .I(pwmWriteZ0Z_0));
    LocalMux I__2037 (
            .O(N__16859),
            .I(pwmWriteZ0Z_0));
    InMux I__2036 (
            .O(N__16854),
            .I(N__16850));
    InMux I__2035 (
            .O(N__16853),
            .I(N__16847));
    LocalMux I__2034 (
            .O(N__16850),
            .I(\QuadInstance7.delayedCh_BZ0Z_1 ));
    LocalMux I__2033 (
            .O(N__16847),
            .I(\QuadInstance7.delayedCh_BZ0Z_1 ));
    InMux I__2032 (
            .O(N__16842),
            .I(N__16836));
    InMux I__2031 (
            .O(N__16841),
            .I(N__16836));
    LocalMux I__2030 (
            .O(N__16836),
            .I(\QuadInstance7.delayedCh_BZ0Z_2 ));
    InMux I__2029 (
            .O(N__16833),
            .I(N__16830));
    LocalMux I__2028 (
            .O(N__16830),
            .I(\PWMInstance1.un1_periodCounter12_1_0_a2_0 ));
    CEMux I__2027 (
            .O(N__16827),
            .I(N__16819));
    CEMux I__2026 (
            .O(N__16826),
            .I(N__16816));
    CEMux I__2025 (
            .O(N__16825),
            .I(N__16813));
    CEMux I__2024 (
            .O(N__16824),
            .I(N__16810));
    CEMux I__2023 (
            .O(N__16823),
            .I(N__16807));
    CEMux I__2022 (
            .O(N__16822),
            .I(N__16804));
    LocalMux I__2021 (
            .O(N__16819),
            .I(N__16800));
    LocalMux I__2020 (
            .O(N__16816),
            .I(N__16795));
    LocalMux I__2019 (
            .O(N__16813),
            .I(N__16795));
    LocalMux I__2018 (
            .O(N__16810),
            .I(N__16792));
    LocalMux I__2017 (
            .O(N__16807),
            .I(N__16789));
    LocalMux I__2016 (
            .O(N__16804),
            .I(N__16786));
    CEMux I__2015 (
            .O(N__16803),
            .I(N__16783));
    Span4Mux_s3_v I__2014 (
            .O(N__16800),
            .I(N__16778));
    Span4Mux_h I__2013 (
            .O(N__16795),
            .I(N__16778));
    Span4Mux_v I__2012 (
            .O(N__16792),
            .I(N__16775));
    Span4Mux_s2_v I__2011 (
            .O(N__16789),
            .I(N__16768));
    Span4Mux_h I__2010 (
            .O(N__16786),
            .I(N__16768));
    LocalMux I__2009 (
            .O(N__16783),
            .I(N__16768));
    Span4Mux_v I__2008 (
            .O(N__16778),
            .I(N__16765));
    Span4Mux_h I__2007 (
            .O(N__16775),
            .I(N__16760));
    Span4Mux_v I__2006 (
            .O(N__16768),
            .I(N__16760));
    Odrv4 I__2005 (
            .O(N__16765),
            .I(\PWMInstance1.pwmWrite_0_1 ));
    Odrv4 I__2004 (
            .O(N__16760),
            .I(\PWMInstance1.pwmWrite_0_1 ));
    InMux I__2003 (
            .O(N__16755),
            .I(N__16746));
    InMux I__2002 (
            .O(N__16754),
            .I(N__16746));
    InMux I__2001 (
            .O(N__16753),
            .I(N__16746));
    LocalMux I__2000 (
            .O(N__16746),
            .I(pwmWriteZ0Z_1));
    CascadeMux I__1999 (
            .O(N__16743),
            .I(N__16739));
    CascadeMux I__1998 (
            .O(N__16742),
            .I(N__16736));
    InMux I__1997 (
            .O(N__16739),
            .I(N__16725));
    InMux I__1996 (
            .O(N__16736),
            .I(N__16725));
    InMux I__1995 (
            .O(N__16735),
            .I(N__16725));
    InMux I__1994 (
            .O(N__16734),
            .I(N__16725));
    LocalMux I__1993 (
            .O(N__16725),
            .I(\PWMInstance1.clkCountZ0Z_1 ));
    InMux I__1992 (
            .O(N__16722),
            .I(N__16710));
    InMux I__1991 (
            .O(N__16721),
            .I(N__16710));
    InMux I__1990 (
            .O(N__16720),
            .I(N__16710));
    InMux I__1989 (
            .O(N__16719),
            .I(N__16710));
    LocalMux I__1988 (
            .O(N__16710),
            .I(\PWMInstance1.clkCountZ0Z_0 ));
    CascadeMux I__1987 (
            .O(N__16707),
            .I(N__16704));
    InMux I__1986 (
            .O(N__16704),
            .I(N__16697));
    InMux I__1985 (
            .O(N__16703),
            .I(N__16697));
    InMux I__1984 (
            .O(N__16702),
            .I(N__16694));
    LocalMux I__1983 (
            .O(N__16697),
            .I(N__16691));
    LocalMux I__1982 (
            .O(N__16694),
            .I(\PWMInstance1.periodCounterZ0Z_16 ));
    Odrv12 I__1981 (
            .O(N__16691),
            .I(\PWMInstance1.periodCounterZ0Z_16 ));
    InMux I__1980 (
            .O(N__16686),
            .I(N__16683));
    LocalMux I__1979 (
            .O(N__16683),
            .I(N__16679));
    InMux I__1978 (
            .O(N__16682),
            .I(N__16675));
    Span4Mux_v I__1977 (
            .O(N__16679),
            .I(N__16672));
    InMux I__1976 (
            .O(N__16678),
            .I(N__16669));
    LocalMux I__1975 (
            .O(N__16675),
            .I(N__16664));
    Span4Mux_v I__1974 (
            .O(N__16672),
            .I(N__16664));
    LocalMux I__1973 (
            .O(N__16669),
            .I(\PWMInstance1.periodCounterZ0Z_7 ));
    Odrv4 I__1972 (
            .O(N__16664),
            .I(\PWMInstance1.periodCounterZ0Z_7 ));
    CascadeMux I__1971 (
            .O(N__16659),
            .I(N__16656));
    InMux I__1970 (
            .O(N__16656),
            .I(N__16652));
    InMux I__1969 (
            .O(N__16655),
            .I(N__16649));
    LocalMux I__1968 (
            .O(N__16652),
            .I(N__16645));
    LocalMux I__1967 (
            .O(N__16649),
            .I(N__16642));
    InMux I__1966 (
            .O(N__16648),
            .I(N__16639));
    Span4Mux_h I__1965 (
            .O(N__16645),
            .I(N__16636));
    Span12Mux_s11_v I__1964 (
            .O(N__16642),
            .I(N__16633));
    LocalMux I__1963 (
            .O(N__16639),
            .I(\PWMInstance1.periodCounterZ0Z_15 ));
    Odrv4 I__1962 (
            .O(N__16636),
            .I(\PWMInstance1.periodCounterZ0Z_15 ));
    Odrv12 I__1961 (
            .O(N__16633),
            .I(\PWMInstance1.periodCounterZ0Z_15 ));
    InMux I__1960 (
            .O(N__16626),
            .I(N__16623));
    LocalMux I__1959 (
            .O(N__16623),
            .I(N__16620));
    Span4Mux_v I__1958 (
            .O(N__16620),
            .I(N__16615));
    InMux I__1957 (
            .O(N__16619),
            .I(N__16612));
    InMux I__1956 (
            .O(N__16618),
            .I(N__16609));
    Span4Mux_v I__1955 (
            .O(N__16615),
            .I(N__16604));
    LocalMux I__1954 (
            .O(N__16612),
            .I(N__16604));
    LocalMux I__1953 (
            .O(N__16609),
            .I(\PWMInstance1.periodCounterZ0Z_1 ));
    Odrv4 I__1952 (
            .O(N__16604),
            .I(\PWMInstance1.periodCounterZ0Z_1 ));
    CascadeMux I__1951 (
            .O(N__16599),
            .I(\PWMInstance1.un1_periodCounter12_1_0_a2_0_6_cascade_ ));
    CascadeMux I__1950 (
            .O(N__16596),
            .I(N__16592));
    InMux I__1949 (
            .O(N__16595),
            .I(N__16589));
    InMux I__1948 (
            .O(N__16592),
            .I(N__16586));
    LocalMux I__1947 (
            .O(N__16589),
            .I(N__16581));
    LocalMux I__1946 (
            .O(N__16586),
            .I(N__16581));
    Span12Mux_s2_v I__1945 (
            .O(N__16581),
            .I(N__16577));
    InMux I__1944 (
            .O(N__16580),
            .I(N__16574));
    Odrv12 I__1943 (
            .O(N__16577),
            .I(\PWMInstance1.periodCounter12 ));
    LocalMux I__1942 (
            .O(N__16574),
            .I(\PWMInstance1.periodCounter12 ));
    InMux I__1941 (
            .O(N__16569),
            .I(N__16566));
    LocalMux I__1940 (
            .O(N__16566),
            .I(N__16563));
    Span4Mux_v I__1939 (
            .O(N__16563),
            .I(N__16560));
    Span4Mux_v I__1938 (
            .O(N__16560),
            .I(N__16557));
    Odrv4 I__1937 (
            .O(N__16557),
            .I(\PWMInstance1.un1_periodCounter12_1_0_a2_0_10 ));
    InMux I__1936 (
            .O(N__16554),
            .I(N__16551));
    LocalMux I__1935 (
            .O(N__16551),
            .I(N__16548));
    Span12Mux_h I__1934 (
            .O(N__16548),
            .I(N__16545));
    Odrv12 I__1933 (
            .O(N__16545),
            .I(\PWMInstance1.un1_periodCounter12_1_0_a2_0_9 ));
    CascadeMux I__1932 (
            .O(N__16542),
            .I(\PWMInstance1.un1_periodCounter12_1_0_a2_0_14_cascade_ ));
    InMux I__1931 (
            .O(N__16539),
            .I(N__16536));
    LocalMux I__1930 (
            .O(N__16536),
            .I(N__16533));
    Span4Mux_v I__1929 (
            .O(N__16533),
            .I(N__16530));
    Span4Mux_v I__1928 (
            .O(N__16530),
            .I(N__16527));
    Odrv4 I__1927 (
            .O(N__16527),
            .I(\PWMInstance1.un1_periodCounter12_1_0_a2_0_12 ));
    CascadeMux I__1926 (
            .O(N__16524),
            .I(N__16518));
    CascadeMux I__1925 (
            .O(N__16523),
            .I(N__16515));
    InMux I__1924 (
            .O(N__16522),
            .I(N__16502));
    InMux I__1923 (
            .O(N__16521),
            .I(N__16495));
    InMux I__1922 (
            .O(N__16518),
            .I(N__16495));
    InMux I__1921 (
            .O(N__16515),
            .I(N__16495));
    InMux I__1920 (
            .O(N__16514),
            .I(N__16484));
    InMux I__1919 (
            .O(N__16513),
            .I(N__16484));
    InMux I__1918 (
            .O(N__16512),
            .I(N__16484));
    InMux I__1917 (
            .O(N__16511),
            .I(N__16484));
    InMux I__1916 (
            .O(N__16510),
            .I(N__16484));
    InMux I__1915 (
            .O(N__16509),
            .I(N__16473));
    InMux I__1914 (
            .O(N__16508),
            .I(N__16473));
    InMux I__1913 (
            .O(N__16507),
            .I(N__16473));
    InMux I__1912 (
            .O(N__16506),
            .I(N__16473));
    InMux I__1911 (
            .O(N__16505),
            .I(N__16473));
    LocalMux I__1910 (
            .O(N__16502),
            .I(\QuadInstance7.un1_count_enable_i_a2_0_1 ));
    LocalMux I__1909 (
            .O(N__16495),
            .I(\QuadInstance7.un1_count_enable_i_a2_0_1 ));
    LocalMux I__1908 (
            .O(N__16484),
            .I(\QuadInstance7.un1_count_enable_i_a2_0_1 ));
    LocalMux I__1907 (
            .O(N__16473),
            .I(\QuadInstance7.un1_count_enable_i_a2_0_1 ));
    InMux I__1906 (
            .O(N__16464),
            .I(N__16459));
    InMux I__1905 (
            .O(N__16463),
            .I(N__16454));
    InMux I__1904 (
            .O(N__16462),
            .I(N__16454));
    LocalMux I__1903 (
            .O(N__16459),
            .I(\QuadInstance7.delayedCh_AZ0Z_1 ));
    LocalMux I__1902 (
            .O(N__16454),
            .I(\QuadInstance7.delayedCh_AZ0Z_1 ));
    CascadeMux I__1901 (
            .O(N__16449),
            .I(N__16446));
    InMux I__1900 (
            .O(N__16446),
            .I(N__16443));
    LocalMux I__1899 (
            .O(N__16443),
            .I(\QuadInstance7.delayedCh_AZ0Z_2 ));
    CascadeMux I__1898 (
            .O(N__16440),
            .I(\QuadInstance7.un1_count_enable_i_a2_0_1_cascade_ ));
    CascadeMux I__1897 (
            .O(N__16437),
            .I(\QuadInstance7.count_enable_cascade_ ));
    InMux I__1896 (
            .O(N__16434),
            .I(N__16431));
    LocalMux I__1895 (
            .O(N__16431),
            .I(\QuadInstance2.Quad_RNO_0_2_10 ));
    InMux I__1894 (
            .O(N__16428),
            .I(N__16425));
    LocalMux I__1893 (
            .O(N__16425),
            .I(\QuadInstance2.Quad_RNO_0_2_14 ));
    InMux I__1892 (
            .O(N__16422),
            .I(N__16419));
    LocalMux I__1891 (
            .O(N__16419),
            .I(\QuadInstance2.Quad_RNO_0_2_12 ));
    InMux I__1890 (
            .O(N__16416),
            .I(N__16413));
    LocalMux I__1889 (
            .O(N__16413),
            .I(N__16410));
    Span12Mux_h I__1888 (
            .O(N__16410),
            .I(N__16407));
    Odrv12 I__1887 (
            .O(N__16407),
            .I(\PWMInstance5.un1_PWMPulseWidthCount_0_I_45_c_RNO_4 ));
    InMux I__1886 (
            .O(N__16404),
            .I(bfn_8_5_0_));
    IoInMux I__1885 (
            .O(N__16401),
            .I(N__16398));
    LocalMux I__1884 (
            .O(N__16398),
            .I(N__16395));
    Span4Mux_s3_v I__1883 (
            .O(N__16395),
            .I(N__16392));
    Sp12to4 I__1882 (
            .O(N__16392),
            .I(N__16389));
    Span12Mux_h I__1881 (
            .O(N__16389),
            .I(N__16386));
    Span12Mux_v I__1880 (
            .O(N__16386),
            .I(N__16382));
    InMux I__1879 (
            .O(N__16385),
            .I(N__16379));
    Odrv12 I__1878 (
            .O(N__16382),
            .I(PWM5_c));
    LocalMux I__1877 (
            .O(N__16379),
            .I(PWM5_c));
    CascadeMux I__1876 (
            .O(N__16374),
            .I(N__16371));
    InMux I__1875 (
            .O(N__16371),
            .I(N__16368));
    LocalMux I__1874 (
            .O(N__16368),
            .I(\PWMInstance1.PWMPulseWidthCountZ0Z_12 ));
    InMux I__1873 (
            .O(N__16365),
            .I(N__16362));
    LocalMux I__1872 (
            .O(N__16362),
            .I(\PWMInstance1.PWMPulseWidthCountZ0Z_10 ));
    CascadeMux I__1871 (
            .O(N__16359),
            .I(N__16356));
    InMux I__1870 (
            .O(N__16356),
            .I(N__16353));
    LocalMux I__1869 (
            .O(N__16353),
            .I(\QuadInstance2.Quad_RNO_0_2_9 ));
    InMux I__1868 (
            .O(N__16350),
            .I(N__16345));
    CascadeMux I__1867 (
            .O(N__16349),
            .I(N__16342));
    InMux I__1866 (
            .O(N__16348),
            .I(N__16339));
    LocalMux I__1865 (
            .O(N__16345),
            .I(N__16336));
    InMux I__1864 (
            .O(N__16342),
            .I(N__16333));
    LocalMux I__1863 (
            .O(N__16339),
            .I(\PWMInstance1.periodCounterZ0Z_11 ));
    Odrv4 I__1862 (
            .O(N__16336),
            .I(\PWMInstance1.periodCounterZ0Z_11 ));
    LocalMux I__1861 (
            .O(N__16333),
            .I(\PWMInstance1.periodCounterZ0Z_11 ));
    InMux I__1860 (
            .O(N__16326),
            .I(\PWMInstance1.un1_periodCounter_2_cry_10 ));
    InMux I__1859 (
            .O(N__16323),
            .I(N__16319));
    InMux I__1858 (
            .O(N__16322),
            .I(N__16315));
    LocalMux I__1857 (
            .O(N__16319),
            .I(N__16312));
    InMux I__1856 (
            .O(N__16318),
            .I(N__16309));
    LocalMux I__1855 (
            .O(N__16315),
            .I(\PWMInstance1.periodCounterZ0Z_12 ));
    Odrv4 I__1854 (
            .O(N__16312),
            .I(\PWMInstance1.periodCounterZ0Z_12 ));
    LocalMux I__1853 (
            .O(N__16309),
            .I(\PWMInstance1.periodCounterZ0Z_12 ));
    InMux I__1852 (
            .O(N__16302),
            .I(\PWMInstance1.un1_periodCounter_2_cry_11 ));
    InMux I__1851 (
            .O(N__16299),
            .I(N__16296));
    LocalMux I__1850 (
            .O(N__16296),
            .I(N__16291));
    InMux I__1849 (
            .O(N__16295),
            .I(N__16288));
    InMux I__1848 (
            .O(N__16294),
            .I(N__16285));
    Span4Mux_h I__1847 (
            .O(N__16291),
            .I(N__16280));
    LocalMux I__1846 (
            .O(N__16288),
            .I(N__16280));
    LocalMux I__1845 (
            .O(N__16285),
            .I(\PWMInstance1.periodCounterZ0Z_13 ));
    Odrv4 I__1844 (
            .O(N__16280),
            .I(\PWMInstance1.periodCounterZ0Z_13 ));
    InMux I__1843 (
            .O(N__16275),
            .I(\PWMInstance1.un1_periodCounter_2_cry_12 ));
    InMux I__1842 (
            .O(N__16272),
            .I(N__16268));
    InMux I__1841 (
            .O(N__16271),
            .I(N__16264));
    LocalMux I__1840 (
            .O(N__16268),
            .I(N__16261));
    InMux I__1839 (
            .O(N__16267),
            .I(N__16258));
    LocalMux I__1838 (
            .O(N__16264),
            .I(\PWMInstance1.periodCounterZ0Z_14 ));
    Odrv4 I__1837 (
            .O(N__16261),
            .I(\PWMInstance1.periodCounterZ0Z_14 ));
    LocalMux I__1836 (
            .O(N__16258),
            .I(\PWMInstance1.periodCounterZ0Z_14 ));
    InMux I__1835 (
            .O(N__16251),
            .I(\PWMInstance1.un1_periodCounter_2_cry_13 ));
    InMux I__1834 (
            .O(N__16248),
            .I(\PWMInstance1.un1_periodCounter_2_cry_14 ));
    InMux I__1833 (
            .O(N__16245),
            .I(bfn_8_3_0_));
    CascadeMux I__1832 (
            .O(N__16242),
            .I(N__16237));
    InMux I__1831 (
            .O(N__16241),
            .I(N__16234));
    InMux I__1830 (
            .O(N__16240),
            .I(N__16229));
    InMux I__1829 (
            .O(N__16237),
            .I(N__16229));
    LocalMux I__1828 (
            .O(N__16234),
            .I(\PWMInstance1.periodCounterZ0Z_3 ));
    LocalMux I__1827 (
            .O(N__16229),
            .I(\PWMInstance1.periodCounterZ0Z_3 ));
    InMux I__1826 (
            .O(N__16224),
            .I(\PWMInstance1.un1_periodCounter_2_cry_2 ));
    InMux I__1825 (
            .O(N__16221),
            .I(N__16216));
    InMux I__1824 (
            .O(N__16220),
            .I(N__16211));
    InMux I__1823 (
            .O(N__16219),
            .I(N__16211));
    LocalMux I__1822 (
            .O(N__16216),
            .I(\PWMInstance1.periodCounterZ0Z_4 ));
    LocalMux I__1821 (
            .O(N__16211),
            .I(\PWMInstance1.periodCounterZ0Z_4 ));
    InMux I__1820 (
            .O(N__16206),
            .I(\PWMInstance1.un1_periodCounter_2_cry_3 ));
    CascadeMux I__1819 (
            .O(N__16203),
            .I(N__16198));
    InMux I__1818 (
            .O(N__16202),
            .I(N__16195));
    InMux I__1817 (
            .O(N__16201),
            .I(N__16190));
    InMux I__1816 (
            .O(N__16198),
            .I(N__16190));
    LocalMux I__1815 (
            .O(N__16195),
            .I(\PWMInstance1.periodCounterZ0Z_5 ));
    LocalMux I__1814 (
            .O(N__16190),
            .I(\PWMInstance1.periodCounterZ0Z_5 ));
    InMux I__1813 (
            .O(N__16185),
            .I(\PWMInstance1.un1_periodCounter_2_cry_4 ));
    CascadeMux I__1812 (
            .O(N__16182),
            .I(N__16179));
    InMux I__1811 (
            .O(N__16179),
            .I(N__16173));
    InMux I__1810 (
            .O(N__16178),
            .I(N__16173));
    LocalMux I__1809 (
            .O(N__16173),
            .I(N__16169));
    InMux I__1808 (
            .O(N__16172),
            .I(N__16166));
    Span4Mux_h I__1807 (
            .O(N__16169),
            .I(N__16163));
    LocalMux I__1806 (
            .O(N__16166),
            .I(\PWMInstance1.periodCounterZ0Z_6 ));
    Odrv4 I__1805 (
            .O(N__16163),
            .I(\PWMInstance1.periodCounterZ0Z_6 ));
    InMux I__1804 (
            .O(N__16158),
            .I(\PWMInstance1.un1_periodCounter_2_cry_5 ));
    InMux I__1803 (
            .O(N__16155),
            .I(\PWMInstance1.un1_periodCounter_2_cry_6 ));
    InMux I__1802 (
            .O(N__16152),
            .I(N__16147));
    InMux I__1801 (
            .O(N__16151),
            .I(N__16144));
    InMux I__1800 (
            .O(N__16150),
            .I(N__16141));
    LocalMux I__1799 (
            .O(N__16147),
            .I(\PWMInstance1.periodCounterZ0Z_8 ));
    LocalMux I__1798 (
            .O(N__16144),
            .I(\PWMInstance1.periodCounterZ0Z_8 ));
    LocalMux I__1797 (
            .O(N__16141),
            .I(\PWMInstance1.periodCounterZ0Z_8 ));
    InMux I__1796 (
            .O(N__16134),
            .I(bfn_8_2_0_));
    CascadeMux I__1795 (
            .O(N__16131),
            .I(N__16126));
    InMux I__1794 (
            .O(N__16130),
            .I(N__16123));
    InMux I__1793 (
            .O(N__16129),
            .I(N__16120));
    InMux I__1792 (
            .O(N__16126),
            .I(N__16117));
    LocalMux I__1791 (
            .O(N__16123),
            .I(\PWMInstance1.periodCounterZ0Z_9 ));
    LocalMux I__1790 (
            .O(N__16120),
            .I(\PWMInstance1.periodCounterZ0Z_9 ));
    LocalMux I__1789 (
            .O(N__16117),
            .I(\PWMInstance1.periodCounterZ0Z_9 ));
    InMux I__1788 (
            .O(N__16110),
            .I(\PWMInstance1.un1_periodCounter_2_cry_8 ));
    InMux I__1787 (
            .O(N__16107),
            .I(N__16104));
    LocalMux I__1786 (
            .O(N__16104),
            .I(N__16099));
    InMux I__1785 (
            .O(N__16103),
            .I(N__16096));
    InMux I__1784 (
            .O(N__16102),
            .I(N__16093));
    Span4Mux_h I__1783 (
            .O(N__16099),
            .I(N__16090));
    LocalMux I__1782 (
            .O(N__16096),
            .I(\PWMInstance1.periodCounterZ0Z_10 ));
    LocalMux I__1781 (
            .O(N__16093),
            .I(\PWMInstance1.periodCounterZ0Z_10 ));
    Odrv4 I__1780 (
            .O(N__16090),
            .I(\PWMInstance1.periodCounterZ0Z_10 ));
    InMux I__1779 (
            .O(N__16083),
            .I(\PWMInstance1.un1_periodCounter_2_cry_9 ));
    InMux I__1778 (
            .O(N__16080),
            .I(\PWMInstance0.un1_periodCounter_2_cry_10 ));
    InMux I__1777 (
            .O(N__16077),
            .I(\PWMInstance0.un1_periodCounter_2_cry_11 ));
    InMux I__1776 (
            .O(N__16074),
            .I(\PWMInstance0.un1_periodCounter_2_cry_12 ));
    InMux I__1775 (
            .O(N__16071),
            .I(\PWMInstance0.un1_periodCounter_2_cry_13 ));
    InMux I__1774 (
            .O(N__16068),
            .I(\PWMInstance0.un1_periodCounter_2_cry_14 ));
    InMux I__1773 (
            .O(N__16065),
            .I(bfn_7_18_0_));
    InMux I__1772 (
            .O(N__16062),
            .I(N__16055));
    InMux I__1771 (
            .O(N__16061),
            .I(N__16055));
    InMux I__1770 (
            .O(N__16060),
            .I(N__16052));
    LocalMux I__1769 (
            .O(N__16055),
            .I(N__16049));
    LocalMux I__1768 (
            .O(N__16052),
            .I(\PWMInstance0.periodCounterZ0Z_16 ));
    Odrv4 I__1767 (
            .O(N__16049),
            .I(\PWMInstance0.periodCounterZ0Z_16 ));
    InMux I__1766 (
            .O(N__16044),
            .I(N__16037));
    InMux I__1765 (
            .O(N__16043),
            .I(N__16037));
    InMux I__1764 (
            .O(N__16042),
            .I(N__16034));
    LocalMux I__1763 (
            .O(N__16037),
            .I(N__16031));
    LocalMux I__1762 (
            .O(N__16034),
            .I(\PWMInstance1.periodCounterZ0Z_0 ));
    Odrv4 I__1761 (
            .O(N__16031),
            .I(\PWMInstance1.periodCounterZ0Z_0 ));
    InMux I__1760 (
            .O(N__16026),
            .I(\PWMInstance1.un1_periodCounter_2_cry_0 ));
    InMux I__1759 (
            .O(N__16023),
            .I(N__16018));
    InMux I__1758 (
            .O(N__16022),
            .I(N__16013));
    InMux I__1757 (
            .O(N__16021),
            .I(N__16013));
    LocalMux I__1756 (
            .O(N__16018),
            .I(\PWMInstance1.periodCounterZ0Z_2 ));
    LocalMux I__1755 (
            .O(N__16013),
            .I(\PWMInstance1.periodCounterZ0Z_2 ));
    InMux I__1754 (
            .O(N__16008),
            .I(\PWMInstance1.un1_periodCounter_2_cry_1 ));
    InMux I__1753 (
            .O(N__16005),
            .I(N__15998));
    InMux I__1752 (
            .O(N__16004),
            .I(N__15998));
    InMux I__1751 (
            .O(N__16003),
            .I(N__15995));
    LocalMux I__1750 (
            .O(N__15998),
            .I(N__15992));
    LocalMux I__1749 (
            .O(N__15995),
            .I(\PWMInstance0.periodCounterZ0Z_2 ));
    Odrv4 I__1748 (
            .O(N__15992),
            .I(\PWMInstance0.periodCounterZ0Z_2 ));
    InMux I__1747 (
            .O(N__15987),
            .I(\PWMInstance0.un1_periodCounter_2_cry_1 ));
    CascadeMux I__1746 (
            .O(N__15984),
            .I(N__15980));
    InMux I__1745 (
            .O(N__15983),
            .I(N__15974));
    InMux I__1744 (
            .O(N__15980),
            .I(N__15974));
    InMux I__1743 (
            .O(N__15979),
            .I(N__15971));
    LocalMux I__1742 (
            .O(N__15974),
            .I(N__15968));
    LocalMux I__1741 (
            .O(N__15971),
            .I(\PWMInstance0.periodCounterZ0Z_3 ));
    Odrv4 I__1740 (
            .O(N__15968),
            .I(\PWMInstance0.periodCounterZ0Z_3 ));
    InMux I__1739 (
            .O(N__15963),
            .I(\PWMInstance0.un1_periodCounter_2_cry_2 ));
    InMux I__1738 (
            .O(N__15960),
            .I(N__15953));
    InMux I__1737 (
            .O(N__15959),
            .I(N__15953));
    InMux I__1736 (
            .O(N__15958),
            .I(N__15950));
    LocalMux I__1735 (
            .O(N__15953),
            .I(N__15947));
    LocalMux I__1734 (
            .O(N__15950),
            .I(\PWMInstance0.periodCounterZ0Z_4 ));
    Odrv4 I__1733 (
            .O(N__15947),
            .I(\PWMInstance0.periodCounterZ0Z_4 ));
    InMux I__1732 (
            .O(N__15942),
            .I(\PWMInstance0.un1_periodCounter_2_cry_3 ));
    CascadeMux I__1731 (
            .O(N__15939),
            .I(N__15935));
    InMux I__1730 (
            .O(N__15938),
            .I(N__15929));
    InMux I__1729 (
            .O(N__15935),
            .I(N__15929));
    InMux I__1728 (
            .O(N__15934),
            .I(N__15926));
    LocalMux I__1727 (
            .O(N__15929),
            .I(N__15923));
    LocalMux I__1726 (
            .O(N__15926),
            .I(\PWMInstance0.periodCounterZ0Z_5 ));
    Odrv4 I__1725 (
            .O(N__15923),
            .I(\PWMInstance0.periodCounterZ0Z_5 ));
    InMux I__1724 (
            .O(N__15918),
            .I(\PWMInstance0.un1_periodCounter_2_cry_4 ));
    InMux I__1723 (
            .O(N__15915),
            .I(\PWMInstance0.un1_periodCounter_2_cry_5 ));
    InMux I__1722 (
            .O(N__15912),
            .I(\PWMInstance0.un1_periodCounter_2_cry_6 ));
    InMux I__1721 (
            .O(N__15909),
            .I(bfn_7_17_0_));
    InMux I__1720 (
            .O(N__15906),
            .I(\PWMInstance0.un1_periodCounter_2_cry_8 ));
    InMux I__1719 (
            .O(N__15903),
            .I(\PWMInstance0.un1_periodCounter_2_cry_9 ));
    InMux I__1718 (
            .O(N__15900),
            .I(N__15894));
    InMux I__1717 (
            .O(N__15899),
            .I(N__15894));
    LocalMux I__1716 (
            .O(N__15894),
            .I(N__15891));
    Odrv12 I__1715 (
            .O(N__15891),
            .I(pwmWrite_fastZ0Z_0));
    CascadeMux I__1714 (
            .O(N__15888),
            .I(N__15883));
    InMux I__1713 (
            .O(N__15887),
            .I(N__15873));
    InMux I__1712 (
            .O(N__15886),
            .I(N__15873));
    InMux I__1711 (
            .O(N__15883),
            .I(N__15873));
    InMux I__1710 (
            .O(N__15882),
            .I(N__15873));
    LocalMux I__1709 (
            .O(N__15873),
            .I(\PWMInstance0.clkCountZ0Z_1 ));
    InMux I__1708 (
            .O(N__15870),
            .I(N__15858));
    InMux I__1707 (
            .O(N__15869),
            .I(N__15858));
    InMux I__1706 (
            .O(N__15868),
            .I(N__15858));
    InMux I__1705 (
            .O(N__15867),
            .I(N__15858));
    LocalMux I__1704 (
            .O(N__15858),
            .I(\PWMInstance0.clkCountZ0Z_0 ));
    CascadeMux I__1703 (
            .O(N__15855),
            .I(\PWMInstance0.periodCounter12_cascade_ ));
    InMux I__1702 (
            .O(N__15852),
            .I(N__15849));
    LocalMux I__1701 (
            .O(N__15849),
            .I(\PWMInstance0.un1_periodCounter12_1_0_a2_0_6 ));
    InMux I__1700 (
            .O(N__15846),
            .I(N__15843));
    LocalMux I__1699 (
            .O(N__15843),
            .I(\PWMInstance0.un1_periodCounter12_1_0_a2_0_10 ));
    CascadeMux I__1698 (
            .O(N__15840),
            .I(\PWMInstance0.un1_periodCounter12_1_0_a2_0_14_cascade_ ));
    InMux I__1697 (
            .O(N__15837),
            .I(N__15834));
    LocalMux I__1696 (
            .O(N__15834),
            .I(\PWMInstance0.un1_periodCounter12_1_0_a2_0_12 ));
    CascadeMux I__1695 (
            .O(N__15831),
            .I(N__15827));
    InMux I__1694 (
            .O(N__15830),
            .I(N__15824));
    InMux I__1693 (
            .O(N__15827),
            .I(N__15821));
    LocalMux I__1692 (
            .O(N__15824),
            .I(\PWMInstance0.periodCounter12 ));
    LocalMux I__1691 (
            .O(N__15821),
            .I(\PWMInstance0.periodCounter12 ));
    InMux I__1690 (
            .O(N__15816),
            .I(\PWMInstance0.un1_periodCounter_2_cry_0 ));
    InMux I__1689 (
            .O(N__15813),
            .I(N__15810));
    LocalMux I__1688 (
            .O(N__15810),
            .I(\PWMInstance0.PWMPulseWidthCountZ0Z_2 ));
    InMux I__1687 (
            .O(N__15807),
            .I(N__15804));
    LocalMux I__1686 (
            .O(N__15804),
            .I(N__15801));
    Odrv4 I__1685 (
            .O(N__15801),
            .I(\PWMInstance0.PWMPulseWidthCountZ0Z_3 ));
    CascadeMux I__1684 (
            .O(N__15798),
            .I(\PWMInstance0.un1_periodCounter12_1_0_a2_0_0_cascade_ ));
    InMux I__1683 (
            .O(N__15795),
            .I(N__15792));
    LocalMux I__1682 (
            .O(N__15792),
            .I(\PWMInstance0.PWMPulseWidthCountZ0Z_5 ));
    InMux I__1681 (
            .O(N__15789),
            .I(N__15786));
    LocalMux I__1680 (
            .O(N__15786),
            .I(\PWMInstance0.PWMPulseWidthCountZ0Z_4 ));
    InMux I__1679 (
            .O(N__15783),
            .I(N__15780));
    LocalMux I__1678 (
            .O(N__15780),
            .I(N__15777));
    Sp12to4 I__1677 (
            .O(N__15777),
            .I(N__15774));
    Odrv12 I__1676 (
            .O(N__15774),
            .I(\PWMInstance1.un1_PWMPulseWidthCount_0_I_45_c_RNO_0 ));
    InMux I__1675 (
            .O(N__15771),
            .I(N__15768));
    LocalMux I__1674 (
            .O(N__15768),
            .I(N__15765));
    Span4Mux_v I__1673 (
            .O(N__15765),
            .I(N__15762));
    Odrv4 I__1672 (
            .O(N__15762),
            .I(\PWMInstance1.un1_PWMPulseWidthCount_0_I_33_c_RNO_0 ));
    InMux I__1671 (
            .O(N__15759),
            .I(N__15756));
    LocalMux I__1670 (
            .O(N__15756),
            .I(N__15753));
    Span4Mux_v I__1669 (
            .O(N__15753),
            .I(N__15750));
    Odrv4 I__1668 (
            .O(N__15750),
            .I(\PWMInstance1.un1_PWMPulseWidthCount_0_I_39_c_RNO_0 ));
    InMux I__1667 (
            .O(N__15747),
            .I(N__15744));
    LocalMux I__1666 (
            .O(N__15744),
            .I(N__15741));
    Odrv12 I__1665 (
            .O(N__15741),
            .I(\PWMInstance1.un1_PWMPulseWidthCount_0_I_21_c_RNO_0 ));
    InMux I__1664 (
            .O(N__15738),
            .I(bfn_7_12_0_));
    IoInMux I__1663 (
            .O(N__15735),
            .I(N__15732));
    LocalMux I__1662 (
            .O(N__15732),
            .I(N__15729));
    Span4Mux_s2_v I__1661 (
            .O(N__15729),
            .I(N__15726));
    Span4Mux_v I__1660 (
            .O(N__15726),
            .I(N__15722));
    InMux I__1659 (
            .O(N__15725),
            .I(N__15719));
    Odrv4 I__1658 (
            .O(N__15722),
            .I(PWM1_c));
    LocalMux I__1657 (
            .O(N__15719),
            .I(PWM1_c));
    InMux I__1656 (
            .O(N__15714),
            .I(N__15711));
    LocalMux I__1655 (
            .O(N__15711),
            .I(N__15708));
    Odrv4 I__1654 (
            .O(N__15708),
            .I(\QuadInstance2.Quad_RNIK13G2Z0Z_14 ));
    InMux I__1653 (
            .O(N__15705),
            .I(N__15701));
    InMux I__1652 (
            .O(N__15704),
            .I(N__15698));
    LocalMux I__1651 (
            .O(N__15701),
            .I(\QuadInstance2.delayedCh_BZ0Z_1 ));
    LocalMux I__1650 (
            .O(N__15698),
            .I(\QuadInstance2.delayedCh_BZ0Z_1 ));
    InMux I__1649 (
            .O(N__15693),
            .I(N__15687));
    InMux I__1648 (
            .O(N__15692),
            .I(N__15687));
    LocalMux I__1647 (
            .O(N__15687),
            .I(\QuadInstance2.delayedCh_BZ0Z_2 ));
    InMux I__1646 (
            .O(N__15684),
            .I(N__15681));
    LocalMux I__1645 (
            .O(N__15681),
            .I(N__15678));
    Odrv12 I__1644 (
            .O(N__15678),
            .I(\PWMInstance1.un1_PWMPulseWidthCount_0_I_1_c_RNO_0 ));
    InMux I__1643 (
            .O(N__15675),
            .I(N__15672));
    LocalMux I__1642 (
            .O(N__15672),
            .I(N__15669));
    Odrv12 I__1641 (
            .O(N__15669),
            .I(\PWMInstance1.un1_PWMPulseWidthCount_0_I_9_c_RNO_0 ));
    InMux I__1640 (
            .O(N__15666),
            .I(N__15663));
    LocalMux I__1639 (
            .O(N__15663),
            .I(N__15660));
    Span4Mux_v I__1638 (
            .O(N__15660),
            .I(N__15657));
    Span4Mux_v I__1637 (
            .O(N__15657),
            .I(N__15654));
    Odrv4 I__1636 (
            .O(N__15654),
            .I(\PWMInstance1.un1_PWMPulseWidthCount_0_I_15_c_RNO_0 ));
    InMux I__1635 (
            .O(N__15651),
            .I(N__15648));
    LocalMux I__1634 (
            .O(N__15648),
            .I(N__15645));
    Span12Mux_v I__1633 (
            .O(N__15645),
            .I(N__15642));
    Odrv12 I__1632 (
            .O(N__15642),
            .I(\PWMInstance1.un1_PWMPulseWidthCount_0_I_27_c_RNO_0 ));
    InMux I__1631 (
            .O(N__15639),
            .I(N__15636));
    LocalMux I__1630 (
            .O(N__15636),
            .I(N__15633));
    Odrv4 I__1629 (
            .O(N__15633),
            .I(\QuadInstance2.un1_Quad_axb_15 ));
    CascadeMux I__1628 (
            .O(N__15630),
            .I(\QuadInstance2.count_enable_cascade_ ));
    CascadeMux I__1627 (
            .O(N__15627),
            .I(N__15624));
    InMux I__1626 (
            .O(N__15624),
            .I(N__15621));
    LocalMux I__1625 (
            .O(N__15621),
            .I(N__15618));
    Odrv4 I__1624 (
            .O(N__15618),
            .I(\QuadInstance2.Quad_RNI1MLE2Z0Z_2 ));
    CascadeMux I__1623 (
            .O(N__15615),
            .I(\QuadInstance2.un1_count_enable_i_a2_0_1_cascade_ ));
    CascadeMux I__1622 (
            .O(N__15612),
            .I(N__15609));
    InMux I__1621 (
            .O(N__15609),
            .I(N__15606));
    LocalMux I__1620 (
            .O(N__15606),
            .I(N__15603));
    Odrv4 I__1619 (
            .O(N__15603),
            .I(\QuadInstance2.Quad_RNI2NLE2Z0Z_3 ));
    CascadeMux I__1618 (
            .O(N__15600),
            .I(N__15597));
    InMux I__1617 (
            .O(N__15597),
            .I(N__15594));
    LocalMux I__1616 (
            .O(N__15594),
            .I(N__15591));
    Odrv4 I__1615 (
            .O(N__15591),
            .I(\QuadInstance2.Quad_RNI4PLE2Z0Z_5 ));
    CascadeMux I__1614 (
            .O(N__15588),
            .I(N__15585));
    InMux I__1613 (
            .O(N__15585),
            .I(N__15582));
    LocalMux I__1612 (
            .O(N__15582),
            .I(N__15579));
    Odrv12 I__1611 (
            .O(N__15579),
            .I(\QuadInstance2.Quad_RNI5QLE2Z0Z_6 ));
    CascadeMux I__1610 (
            .O(N__15576),
            .I(N__15571));
    CascadeMux I__1609 (
            .O(N__15575),
            .I(N__15568));
    InMux I__1608 (
            .O(N__15574),
            .I(N__15565));
    InMux I__1607 (
            .O(N__15571),
            .I(N__15560));
    InMux I__1606 (
            .O(N__15568),
            .I(N__15560));
    LocalMux I__1605 (
            .O(N__15565),
            .I(\QuadInstance2.delayedCh_AZ0Z_1 ));
    LocalMux I__1604 (
            .O(N__15560),
            .I(\QuadInstance2.delayedCh_AZ0Z_1 ));
    InMux I__1603 (
            .O(N__15555),
            .I(N__15552));
    LocalMux I__1602 (
            .O(N__15552),
            .I(\QuadInstance2.delayedCh_AZ0Z_2 ));
    InMux I__1601 (
            .O(N__15549),
            .I(\QuadInstance2.un1_Quad_cry_14 ));
    CascadeMux I__1600 (
            .O(N__15546),
            .I(N__15543));
    InMux I__1599 (
            .O(N__15543),
            .I(N__15540));
    LocalMux I__1598 (
            .O(N__15540),
            .I(\QuadInstance2.Quad_RNI8TLE2Z0Z_9 ));
    CascadeMux I__1597 (
            .O(N__15537),
            .I(N__15534));
    InMux I__1596 (
            .O(N__15534),
            .I(N__15531));
    LocalMux I__1595 (
            .O(N__15531),
            .I(\QuadInstance2.Quad_RNIHU2G2Z0Z_11 ));
    CascadeMux I__1594 (
            .O(N__15528),
            .I(N__15525));
    InMux I__1593 (
            .O(N__15525),
            .I(N__15522));
    LocalMux I__1592 (
            .O(N__15522),
            .I(N__15519));
    Odrv4 I__1591 (
            .O(N__15519),
            .I(\QuadInstance2.Quad_RNI0LLE2Z0Z_1 ));
    CascadeMux I__1590 (
            .O(N__15516),
            .I(N__15513));
    InMux I__1589 (
            .O(N__15513),
            .I(N__15510));
    LocalMux I__1588 (
            .O(N__15510),
            .I(\QuadInstance2.Quad_RNIGT2G2Z0Z_10 ));
    CascadeMux I__1587 (
            .O(N__15507),
            .I(N__15504));
    InMux I__1586 (
            .O(N__15504),
            .I(N__15501));
    LocalMux I__1585 (
            .O(N__15501),
            .I(\QuadInstance2.Quad_RNIIV2G2Z0Z_12 ));
    CascadeMux I__1584 (
            .O(N__15498),
            .I(N__15495));
    InMux I__1583 (
            .O(N__15495),
            .I(N__15492));
    LocalMux I__1582 (
            .O(N__15492),
            .I(N__15489));
    Odrv4 I__1581 (
            .O(N__15489),
            .I(\QuadInstance2.Quad_RNI6RLE2Z0Z_7 ));
    CascadeMux I__1580 (
            .O(N__15486),
            .I(N__15483));
    InMux I__1579 (
            .O(N__15483),
            .I(N__15480));
    LocalMux I__1578 (
            .O(N__15480),
            .I(\QuadInstance2.Quad_RNI7SLE2Z0Z_8 ));
    CascadeMux I__1577 (
            .O(N__15477),
            .I(N__15474));
    InMux I__1576 (
            .O(N__15474),
            .I(N__15471));
    LocalMux I__1575 (
            .O(N__15471),
            .I(N__15468));
    Odrv4 I__1574 (
            .O(N__15468),
            .I(\QuadInstance2.Quad_RNI3OLE2Z0Z_4 ));
    InMux I__1573 (
            .O(N__15465),
            .I(\QuadInstance2.un1_Quad_cry_5 ));
    InMux I__1572 (
            .O(N__15462),
            .I(\QuadInstance2.un1_Quad_cry_6 ));
    InMux I__1571 (
            .O(N__15459),
            .I(bfn_7_7_0_));
    InMux I__1570 (
            .O(N__15456),
            .I(\QuadInstance2.un1_Quad_cry_8 ));
    InMux I__1569 (
            .O(N__15453),
            .I(\QuadInstance2.un1_Quad_cry_9 ));
    InMux I__1568 (
            .O(N__15450),
            .I(\QuadInstance2.un1_Quad_cry_10 ));
    InMux I__1567 (
            .O(N__15447),
            .I(\QuadInstance2.un1_Quad_cry_11 ));
    InMux I__1566 (
            .O(N__15444),
            .I(\QuadInstance2.un1_Quad_cry_12 ));
    InMux I__1565 (
            .O(N__15441),
            .I(\QuadInstance2.un1_Quad_cry_13 ));
    InMux I__1564 (
            .O(N__15438),
            .I(N__15435));
    LocalMux I__1563 (
            .O(N__15435),
            .I(\PWMInstance1.PWMPulseWidthCountZ0Z_15 ));
    CascadeMux I__1562 (
            .O(N__15432),
            .I(N__15429));
    InMux I__1561 (
            .O(N__15429),
            .I(N__15426));
    LocalMux I__1560 (
            .O(N__15426),
            .I(N__15423));
    Span4Mux_h I__1559 (
            .O(N__15423),
            .I(N__15420));
    Odrv4 I__1558 (
            .O(N__15420),
            .I(\PWMInstance1.PWMPulseWidthCountZ0Z_11 ));
    InMux I__1557 (
            .O(N__15417),
            .I(N__15414));
    LocalMux I__1556 (
            .O(N__15414),
            .I(\PWMInstance1.PWMPulseWidthCountZ0Z_13 ));
    InMux I__1555 (
            .O(N__15411),
            .I(\QuadInstance2.un1_Quad_cry_0 ));
    InMux I__1554 (
            .O(N__15408),
            .I(\QuadInstance2.un1_Quad_cry_1 ));
    InMux I__1553 (
            .O(N__15405),
            .I(\QuadInstance2.un1_Quad_cry_2 ));
    InMux I__1552 (
            .O(N__15402),
            .I(\QuadInstance2.un1_Quad_cry_3 ));
    InMux I__1551 (
            .O(N__15399),
            .I(\QuadInstance2.un1_Quad_cry_4 ));
    CascadeMux I__1550 (
            .O(N__15396),
            .I(N__15393));
    InMux I__1549 (
            .O(N__15393),
            .I(N__15390));
    LocalMux I__1548 (
            .O(N__15390),
            .I(\PWMInstance1.PWMPulseWidthCountZ0Z_0 ));
    InMux I__1547 (
            .O(N__15387),
            .I(N__15384));
    LocalMux I__1546 (
            .O(N__15384),
            .I(\PWMInstance1.PWMPulseWidthCountZ0Z_1 ));
    CascadeMux I__1545 (
            .O(N__15381),
            .I(N__15378));
    InMux I__1544 (
            .O(N__15378),
            .I(N__15375));
    LocalMux I__1543 (
            .O(N__15375),
            .I(N__15372));
    Span4Mux_s3_v I__1542 (
            .O(N__15372),
            .I(N__15369));
    Odrv4 I__1541 (
            .O(N__15369),
            .I(\PWMInstance1.PWMPulseWidthCountZ0Z_7 ));
    InMux I__1540 (
            .O(N__15366),
            .I(N__15363));
    LocalMux I__1539 (
            .O(N__15363),
            .I(N__15360));
    Span4Mux_s3_v I__1538 (
            .O(N__15360),
            .I(N__15357));
    Odrv4 I__1537 (
            .O(N__15357),
            .I(\PWMInstance1.PWMPulseWidthCountZ0Z_8 ));
    InMux I__1536 (
            .O(N__15354),
            .I(N__15351));
    LocalMux I__1535 (
            .O(N__15351),
            .I(N__15348));
    Odrv4 I__1534 (
            .O(N__15348),
            .I(\PWMInstance1.PWMPulseWidthCountZ0Z_5 ));
    InMux I__1533 (
            .O(N__15345),
            .I(N__15342));
    LocalMux I__1532 (
            .O(N__15342),
            .I(N__15339));
    Odrv4 I__1531 (
            .O(N__15339),
            .I(\PWMInstance1.PWMPulseWidthCountZ0Z_9 ));
    InMux I__1530 (
            .O(N__15336),
            .I(N__15333));
    LocalMux I__1529 (
            .O(N__15333),
            .I(\PWMInstance1.PWMPulseWidthCountZ0Z_6 ));
    InMux I__1528 (
            .O(N__15330),
            .I(N__15327));
    LocalMux I__1527 (
            .O(N__15327),
            .I(N__15324));
    Span4Mux_h I__1526 (
            .O(N__15324),
            .I(N__15321));
    Odrv4 I__1525 (
            .O(N__15321),
            .I(\PWMInstance1.PWMPulseWidthCountZ0Z_14 ));
    InMux I__1524 (
            .O(N__15318),
            .I(N__15315));
    LocalMux I__1523 (
            .O(N__15315),
            .I(\PWMInstance1.PWMPulseWidthCountZ0Z_2 ));
    InMux I__1522 (
            .O(N__15312),
            .I(N__15309));
    LocalMux I__1521 (
            .O(N__15309),
            .I(N__15306));
    Odrv4 I__1520 (
            .O(N__15306),
            .I(\PWMInstance1.PWMPulseWidthCountZ0Z_3 ));
    CascadeMux I__1519 (
            .O(N__15303),
            .I(\PWMInstance1.un1_periodCounter12_1_0_a2_0_0_cascade_ ));
    InMux I__1518 (
            .O(N__15300),
            .I(N__15297));
    LocalMux I__1517 (
            .O(N__15297),
            .I(\PWMInstance1.PWMPulseWidthCountZ0Z_4 ));
    InMux I__1516 (
            .O(N__15294),
            .I(N__15291));
    LocalMux I__1515 (
            .O(N__15291),
            .I(N__15288));
    Odrv4 I__1514 (
            .O(N__15288),
            .I(\PWMInstance7.PWMPulseWidthCountZ0Z_1 ));
    InMux I__1513 (
            .O(N__15285),
            .I(N__15282));
    LocalMux I__1512 (
            .O(N__15282),
            .I(\PWMInstance7.PWMPulseWidthCountZ0Z_0 ));
    CEMux I__1511 (
            .O(N__15279),
            .I(N__15276));
    LocalMux I__1510 (
            .O(N__15276),
            .I(N__15272));
    CEMux I__1509 (
            .O(N__15275),
            .I(N__15267));
    Span4Mux_v I__1508 (
            .O(N__15272),
            .I(N__15263));
    CEMux I__1507 (
            .O(N__15271),
            .I(N__15260));
    CEMux I__1506 (
            .O(N__15270),
            .I(N__15257));
    LocalMux I__1505 (
            .O(N__15267),
            .I(N__15254));
    CEMux I__1504 (
            .O(N__15266),
            .I(N__15251));
    Span4Mux_v I__1503 (
            .O(N__15263),
            .I(N__15246));
    LocalMux I__1502 (
            .O(N__15260),
            .I(N__15246));
    LocalMux I__1501 (
            .O(N__15257),
            .I(N__15243));
    Span4Mux_v I__1500 (
            .O(N__15254),
            .I(N__15240));
    LocalMux I__1499 (
            .O(N__15251),
            .I(N__15237));
    Span4Mux_v I__1498 (
            .O(N__15246),
            .I(N__15232));
    Span4Mux_h I__1497 (
            .O(N__15243),
            .I(N__15232));
    Span4Mux_h I__1496 (
            .O(N__15240),
            .I(N__15229));
    Span4Mux_h I__1495 (
            .O(N__15237),
            .I(N__15226));
    Odrv4 I__1494 (
            .O(N__15232),
            .I(\PWMInstance7.pwmWrite_0_7 ));
    Odrv4 I__1493 (
            .O(N__15229),
            .I(\PWMInstance7.pwmWrite_0_7 ));
    Odrv4 I__1492 (
            .O(N__15226),
            .I(\PWMInstance7.pwmWrite_0_7 ));
    InMux I__1491 (
            .O(N__15219),
            .I(N__15216));
    LocalMux I__1490 (
            .O(N__15216),
            .I(\PWMInstance5.PWMPulseWidthCountZ0Z_9 ));
    InMux I__1489 (
            .O(N__15213),
            .I(N__15210));
    LocalMux I__1488 (
            .O(N__15210),
            .I(\PWMInstance5.PWMPulseWidthCountZ0Z_8 ));
    IoInMux I__1487 (
            .O(N__15207),
            .I(N__15204));
    LocalMux I__1486 (
            .O(N__15204),
            .I(RST_c_i));
    InMux I__1485 (
            .O(N__15201),
            .I(N__15198));
    LocalMux I__1484 (
            .O(N__15198),
            .I(ch0_B_c));
    InMux I__1483 (
            .O(N__15195),
            .I(N__15192));
    LocalMux I__1482 (
            .O(N__15192),
            .I(N__15189));
    Odrv4 I__1481 (
            .O(N__15189),
            .I(\PWMInstance7.PWMPulseWidthCountZ0Z_8 ));
    InMux I__1480 (
            .O(N__15186),
            .I(N__15183));
    LocalMux I__1479 (
            .O(N__15183),
            .I(\PWMInstance7.PWMPulseWidthCountZ0Z_13 ));
    InMux I__1478 (
            .O(N__15180),
            .I(N__15177));
    LocalMux I__1477 (
            .O(N__15177),
            .I(N__15174));
    Odrv4 I__1476 (
            .O(N__15174),
            .I(\PWMInstance7.PWMPulseWidthCountZ0Z_11 ));
    InMux I__1475 (
            .O(N__15171),
            .I(N__15168));
    LocalMux I__1474 (
            .O(N__15168),
            .I(\PWMInstance7.PWMPulseWidthCountZ0Z_12 ));
    InMux I__1473 (
            .O(N__15165),
            .I(N__15162));
    LocalMux I__1472 (
            .O(N__15162),
            .I(N__15159));
    Odrv4 I__1471 (
            .O(N__15159),
            .I(\PWMInstance7.PWMPulseWidthCountZ0Z_5 ));
    InMux I__1470 (
            .O(N__15156),
            .I(N__15153));
    LocalMux I__1469 (
            .O(N__15153),
            .I(N__15150));
    Odrv4 I__1468 (
            .O(N__15150),
            .I(\PWMInstance7.PWMPulseWidthCountZ0Z_4 ));
    CascadeMux I__1467 (
            .O(N__15147),
            .I(N__15144));
    InMux I__1466 (
            .O(N__15144),
            .I(N__15141));
    LocalMux I__1465 (
            .O(N__15141),
            .I(\PWMInstance7.PWMPulseWidthCountZ0Z_7 ));
    InMux I__1464 (
            .O(N__15138),
            .I(N__15135));
    LocalMux I__1463 (
            .O(N__15135),
            .I(N__15132));
    Odrv4 I__1462 (
            .O(N__15132),
            .I(\PWMInstance7.PWMPulseWidthCountZ0Z_6 ));
    CascadeMux I__1461 (
            .O(N__15129),
            .I(N__15126));
    InMux I__1460 (
            .O(N__15126),
            .I(N__15123));
    LocalMux I__1459 (
            .O(N__15123),
            .I(\PWMInstance7.PWMPulseWidthCountZ0Z_15 ));
    InMux I__1458 (
            .O(N__15120),
            .I(N__15115));
    InMux I__1457 (
            .O(N__15119),
            .I(N__15112));
    InMux I__1456 (
            .O(N__15118),
            .I(N__15109));
    LocalMux I__1455 (
            .O(N__15115),
            .I(N__15106));
    LocalMux I__1454 (
            .O(N__15112),
            .I(N__15103));
    LocalMux I__1453 (
            .O(N__15109),
            .I(\PWMInstance7.periodCounterZ0Z_12 ));
    Odrv4 I__1452 (
            .O(N__15106),
            .I(\PWMInstance7.periodCounterZ0Z_12 ));
    Odrv4 I__1451 (
            .O(N__15103),
            .I(\PWMInstance7.periodCounterZ0Z_12 ));
    CascadeMux I__1450 (
            .O(N__15096),
            .I(N__15092));
    CascadeMux I__1449 (
            .O(N__15095),
            .I(N__15089));
    InMux I__1448 (
            .O(N__15092),
            .I(N__15085));
    InMux I__1447 (
            .O(N__15089),
            .I(N__15082));
    InMux I__1446 (
            .O(N__15088),
            .I(N__15079));
    LocalMux I__1445 (
            .O(N__15085),
            .I(N__15074));
    LocalMux I__1444 (
            .O(N__15082),
            .I(N__15074));
    LocalMux I__1443 (
            .O(N__15079),
            .I(\PWMInstance7.periodCounterZ0Z_13 ));
    Odrv4 I__1442 (
            .O(N__15074),
            .I(\PWMInstance7.periodCounterZ0Z_13 ));
    CascadeMux I__1441 (
            .O(N__15069),
            .I(N__15066));
    InMux I__1440 (
            .O(N__15066),
            .I(N__15063));
    LocalMux I__1439 (
            .O(N__15063),
            .I(\PWMInstance7.un1_PWMPulseWidthCount_0_I_39_c_RNO_6 ));
    InMux I__1438 (
            .O(N__15060),
            .I(N__15057));
    LocalMux I__1437 (
            .O(N__15057),
            .I(N__15052));
    InMux I__1436 (
            .O(N__15056),
            .I(N__15049));
    InMux I__1435 (
            .O(N__15055),
            .I(N__15046));
    Span4Mux_h I__1434 (
            .O(N__15052),
            .I(N__15043));
    LocalMux I__1433 (
            .O(N__15049),
            .I(\PWMInstance7.periodCounterZ0Z_0 ));
    LocalMux I__1432 (
            .O(N__15046),
            .I(\PWMInstance7.periodCounterZ0Z_0 ));
    Odrv4 I__1431 (
            .O(N__15043),
            .I(\PWMInstance7.periodCounterZ0Z_0 ));
    CascadeMux I__1430 (
            .O(N__15036),
            .I(N__15033));
    InMux I__1429 (
            .O(N__15033),
            .I(N__15030));
    LocalMux I__1428 (
            .O(N__15030),
            .I(N__15025));
    InMux I__1427 (
            .O(N__15029),
            .I(N__15022));
    InMux I__1426 (
            .O(N__15028),
            .I(N__15019));
    Span4Mux_h I__1425 (
            .O(N__15025),
            .I(N__15016));
    LocalMux I__1424 (
            .O(N__15022),
            .I(\PWMInstance7.periodCounterZ0Z_1 ));
    LocalMux I__1423 (
            .O(N__15019),
            .I(\PWMInstance7.periodCounterZ0Z_1 ));
    Odrv4 I__1422 (
            .O(N__15016),
            .I(\PWMInstance7.periodCounterZ0Z_1 ));
    InMux I__1421 (
            .O(N__15009),
            .I(N__15006));
    LocalMux I__1420 (
            .O(N__15006),
            .I(\PWMInstance7.un1_PWMPulseWidthCount_0_I_1_c_RNO_6 ));
    InMux I__1419 (
            .O(N__15003),
            .I(N__15000));
    LocalMux I__1418 (
            .O(N__15000),
            .I(N__14995));
    InMux I__1417 (
            .O(N__14999),
            .I(N__14992));
    InMux I__1416 (
            .O(N__14998),
            .I(N__14989));
    Span4Mux_h I__1415 (
            .O(N__14995),
            .I(N__14986));
    LocalMux I__1414 (
            .O(N__14992),
            .I(\PWMInstance7.periodCounterZ0Z_6 ));
    LocalMux I__1413 (
            .O(N__14989),
            .I(\PWMInstance7.periodCounterZ0Z_6 ));
    Odrv4 I__1412 (
            .O(N__14986),
            .I(\PWMInstance7.periodCounterZ0Z_6 ));
    InMux I__1411 (
            .O(N__14979),
            .I(N__14976));
    LocalMux I__1410 (
            .O(N__14976),
            .I(N__14972));
    InMux I__1409 (
            .O(N__14975),
            .I(N__14968));
    Span4Mux_h I__1408 (
            .O(N__14972),
            .I(N__14965));
    InMux I__1407 (
            .O(N__14971),
            .I(N__14962));
    LocalMux I__1406 (
            .O(N__14968),
            .I(\PWMInstance7.periodCounterZ0Z_7 ));
    Odrv4 I__1405 (
            .O(N__14965),
            .I(\PWMInstance7.periodCounterZ0Z_7 ));
    LocalMux I__1404 (
            .O(N__14962),
            .I(\PWMInstance7.periodCounterZ0Z_7 ));
    InMux I__1403 (
            .O(N__14955),
            .I(N__14952));
    LocalMux I__1402 (
            .O(N__14952),
            .I(\PWMInstance7.un1_PWMPulseWidthCount_0_I_27_c_RNO_6 ));
    InMux I__1401 (
            .O(N__14949),
            .I(N__14946));
    LocalMux I__1400 (
            .O(N__14946),
            .I(N__14943));
    Odrv12 I__1399 (
            .O(N__14943),
            .I(\PWMInstance7.un1_periodCounter12_1_0_a2_0 ));
    CascadeMux I__1398 (
            .O(N__14940),
            .I(N__14935));
    InMux I__1397 (
            .O(N__14939),
            .I(N__14930));
    InMux I__1396 (
            .O(N__14938),
            .I(N__14930));
    InMux I__1395 (
            .O(N__14935),
            .I(N__14924));
    LocalMux I__1394 (
            .O(N__14930),
            .I(N__14921));
    InMux I__1393 (
            .O(N__14929),
            .I(N__14918));
    InMux I__1392 (
            .O(N__14928),
            .I(N__14915));
    InMux I__1391 (
            .O(N__14927),
            .I(N__14912));
    LocalMux I__1390 (
            .O(N__14924),
            .I(N__14909));
    Odrv4 I__1389 (
            .O(N__14921),
            .I(\PWMInstance7.out_0_sqmuxa ));
    LocalMux I__1388 (
            .O(N__14918),
            .I(\PWMInstance7.out_0_sqmuxa ));
    LocalMux I__1387 (
            .O(N__14915),
            .I(\PWMInstance7.out_0_sqmuxa ));
    LocalMux I__1386 (
            .O(N__14912),
            .I(\PWMInstance7.out_0_sqmuxa ));
    Odrv4 I__1385 (
            .O(N__14909),
            .I(\PWMInstance7.out_0_sqmuxa ));
    InMux I__1384 (
            .O(N__14898),
            .I(bfn_3_11_0_));
    IoInMux I__1383 (
            .O(N__14895),
            .I(N__14892));
    LocalMux I__1382 (
            .O(N__14892),
            .I(N__14889));
    Span4Mux_s3_v I__1381 (
            .O(N__14889),
            .I(N__14886));
    Span4Mux_h I__1380 (
            .O(N__14886),
            .I(N__14883));
    Span4Mux_v I__1379 (
            .O(N__14883),
            .I(N__14879));
    InMux I__1378 (
            .O(N__14882),
            .I(N__14876));
    Odrv4 I__1377 (
            .O(N__14879),
            .I(PWM7_c));
    LocalMux I__1376 (
            .O(N__14876),
            .I(PWM7_c));
    InMux I__1375 (
            .O(N__14871),
            .I(N__14865));
    InMux I__1374 (
            .O(N__14870),
            .I(N__14865));
    LocalMux I__1373 (
            .O(N__14865),
            .I(pwmWrite_fastZ0Z_7));
    InMux I__1372 (
            .O(N__14862),
            .I(N__14859));
    LocalMux I__1371 (
            .O(N__14859),
            .I(\PWMInstance7.PWMPulseWidthCountZ0Z_9 ));
    InMux I__1370 (
            .O(N__14856),
            .I(N__14853));
    LocalMux I__1369 (
            .O(N__14853),
            .I(\PWMInstance7.PWMPulseWidthCountZ0Z_10 ));
    InMux I__1368 (
            .O(N__14850),
            .I(N__14847));
    LocalMux I__1367 (
            .O(N__14847),
            .I(\PWMInstance7.PWMPulseWidthCountZ0Z_3 ));
    InMux I__1366 (
            .O(N__14844),
            .I(N__14839));
    InMux I__1365 (
            .O(N__14843),
            .I(N__14836));
    InMux I__1364 (
            .O(N__14842),
            .I(N__14833));
    LocalMux I__1363 (
            .O(N__14839),
            .I(N__14828));
    LocalMux I__1362 (
            .O(N__14836),
            .I(N__14828));
    LocalMux I__1361 (
            .O(N__14833),
            .I(N__14825));
    Odrv4 I__1360 (
            .O(N__14828),
            .I(\PWMInstance7.periodCounterZ0Z_15 ));
    Odrv4 I__1359 (
            .O(N__14825),
            .I(\PWMInstance7.periodCounterZ0Z_15 ));
    InMux I__1358 (
            .O(N__14820),
            .I(N__14816));
    InMux I__1357 (
            .O(N__14819),
            .I(N__14813));
    LocalMux I__1356 (
            .O(N__14816),
            .I(N__14807));
    LocalMux I__1355 (
            .O(N__14813),
            .I(N__14807));
    InMux I__1354 (
            .O(N__14812),
            .I(N__14804));
    Odrv4 I__1353 (
            .O(N__14807),
            .I(\PWMInstance7.periodCounterZ0Z_14 ));
    LocalMux I__1352 (
            .O(N__14804),
            .I(\PWMInstance7.periodCounterZ0Z_14 ));
    InMux I__1351 (
            .O(N__14799),
            .I(N__14796));
    LocalMux I__1350 (
            .O(N__14796),
            .I(\PWMInstance7.un1_PWMPulseWidthCount_0_I_21_c_RNO_6 ));
    InMux I__1349 (
            .O(N__14793),
            .I(N__14790));
    LocalMux I__1348 (
            .O(N__14790),
            .I(\PWMInstance7.PWMPulseWidthCountZ0Z_14 ));
    InMux I__1347 (
            .O(N__14787),
            .I(N__14782));
    InMux I__1346 (
            .O(N__14786),
            .I(N__14777));
    InMux I__1345 (
            .O(N__14785),
            .I(N__14777));
    LocalMux I__1344 (
            .O(N__14782),
            .I(\PWMInstance7.periodCounterZ0Z_4 ));
    LocalMux I__1343 (
            .O(N__14777),
            .I(\PWMInstance7.periodCounterZ0Z_4 ));
    CascadeMux I__1342 (
            .O(N__14772),
            .I(N__14767));
    InMux I__1341 (
            .O(N__14771),
            .I(N__14764));
    InMux I__1340 (
            .O(N__14770),
            .I(N__14759));
    InMux I__1339 (
            .O(N__14767),
            .I(N__14759));
    LocalMux I__1338 (
            .O(N__14764),
            .I(\PWMInstance7.periodCounterZ0Z_5 ));
    LocalMux I__1337 (
            .O(N__14759),
            .I(\PWMInstance7.periodCounterZ0Z_5 ));
    InMux I__1336 (
            .O(N__14754),
            .I(N__14749));
    InMux I__1335 (
            .O(N__14753),
            .I(N__14744));
    InMux I__1334 (
            .O(N__14752),
            .I(N__14744));
    LocalMux I__1333 (
            .O(N__14749),
            .I(\PWMInstance7.periodCounterZ0Z_8 ));
    LocalMux I__1332 (
            .O(N__14744),
            .I(\PWMInstance7.periodCounterZ0Z_8 ));
    CascadeMux I__1331 (
            .O(N__14739),
            .I(N__14734));
    InMux I__1330 (
            .O(N__14738),
            .I(N__14731));
    InMux I__1329 (
            .O(N__14737),
            .I(N__14726));
    InMux I__1328 (
            .O(N__14734),
            .I(N__14726));
    LocalMux I__1327 (
            .O(N__14731),
            .I(\PWMInstance7.periodCounterZ0Z_9 ));
    LocalMux I__1326 (
            .O(N__14726),
            .I(\PWMInstance7.periodCounterZ0Z_9 ));
    InMux I__1325 (
            .O(N__14721),
            .I(N__14718));
    LocalMux I__1324 (
            .O(N__14718),
            .I(N__14715));
    Odrv12 I__1323 (
            .O(N__14715),
            .I(\PWMInstance7.un1_PWMPulseWidthCount_0_I_9_c_RNO_6 ));
    InMux I__1322 (
            .O(N__14712),
            .I(N__14709));
    LocalMux I__1321 (
            .O(N__14709),
            .I(\PWMInstance7.un1_PWMPulseWidthCount_0_I_15_c_RNO_6 ));
    InMux I__1320 (
            .O(N__14706),
            .I(N__14703));
    LocalMux I__1319 (
            .O(N__14703),
            .I(\PWMInstance7.un1_PWMPulseWidthCount_0_I_45_c_RNO_6 ));
    InMux I__1318 (
            .O(N__14700),
            .I(N__14697));
    LocalMux I__1317 (
            .O(N__14697),
            .I(\PWMInstance7.un1_PWMPulseWidthCount_0_I_33_c_RNO_6 ));
    InMux I__1316 (
            .O(N__14694),
            .I(N__14682));
    InMux I__1315 (
            .O(N__14693),
            .I(N__14682));
    InMux I__1314 (
            .O(N__14692),
            .I(N__14682));
    InMux I__1313 (
            .O(N__14691),
            .I(N__14682));
    LocalMux I__1312 (
            .O(N__14682),
            .I(\PWMInstance7.clkCountZ0Z_0 ));
    CascadeMux I__1311 (
            .O(N__14679),
            .I(N__14675));
    CascadeMux I__1310 (
            .O(N__14678),
            .I(N__14672));
    InMux I__1309 (
            .O(N__14675),
            .I(N__14661));
    InMux I__1308 (
            .O(N__14672),
            .I(N__14661));
    InMux I__1307 (
            .O(N__14671),
            .I(N__14661));
    InMux I__1306 (
            .O(N__14670),
            .I(N__14661));
    LocalMux I__1305 (
            .O(N__14661),
            .I(\PWMInstance7.clkCountZ0Z_1 ));
    InMux I__1304 (
            .O(N__14658),
            .I(N__14655));
    LocalMux I__1303 (
            .O(N__14655),
            .I(\PWMInstance7.PWMPulseWidthCountZ0Z_2 ));
    InMux I__1302 (
            .O(N__14652),
            .I(N__14647));
    InMux I__1301 (
            .O(N__14651),
            .I(N__14642));
    InMux I__1300 (
            .O(N__14650),
            .I(N__14642));
    LocalMux I__1299 (
            .O(N__14647),
            .I(\PWMInstance7.periodCounterZ0Z_2 ));
    LocalMux I__1298 (
            .O(N__14642),
            .I(\PWMInstance7.periodCounterZ0Z_2 ));
    CascadeMux I__1297 (
            .O(N__14637),
            .I(N__14632));
    InMux I__1296 (
            .O(N__14636),
            .I(N__14629));
    InMux I__1295 (
            .O(N__14635),
            .I(N__14626));
    InMux I__1294 (
            .O(N__14632),
            .I(N__14623));
    LocalMux I__1293 (
            .O(N__14629),
            .I(\PWMInstance7.periodCounterZ0Z_3 ));
    LocalMux I__1292 (
            .O(N__14626),
            .I(\PWMInstance7.periodCounterZ0Z_3 ));
    LocalMux I__1291 (
            .O(N__14623),
            .I(\PWMInstance7.periodCounterZ0Z_3 ));
    CascadeMux I__1290 (
            .O(N__14616),
            .I(N__14612));
    InMux I__1289 (
            .O(N__14615),
            .I(N__14608));
    InMux I__1288 (
            .O(N__14612),
            .I(N__14603));
    InMux I__1287 (
            .O(N__14611),
            .I(N__14603));
    LocalMux I__1286 (
            .O(N__14608),
            .I(\PWMInstance7.periodCounterZ0Z_11 ));
    LocalMux I__1285 (
            .O(N__14603),
            .I(\PWMInstance7.periodCounterZ0Z_11 ));
    CascadeMux I__1284 (
            .O(N__14598),
            .I(N__14593));
    CascadeMux I__1283 (
            .O(N__14597),
            .I(N__14590));
    InMux I__1282 (
            .O(N__14596),
            .I(N__14587));
    InMux I__1281 (
            .O(N__14593),
            .I(N__14582));
    InMux I__1280 (
            .O(N__14590),
            .I(N__14582));
    LocalMux I__1279 (
            .O(N__14587),
            .I(\PWMInstance7.periodCounterZ0Z_10 ));
    LocalMux I__1278 (
            .O(N__14582),
            .I(\PWMInstance7.periodCounterZ0Z_10 ));
    InMux I__1277 (
            .O(N__14577),
            .I(N__14574));
    LocalMux I__1276 (
            .O(N__14574),
            .I(\PWMInstance7.un1_periodCounter12_1_0_a2_0_0 ));
    InMux I__1275 (
            .O(N__14571),
            .I(N__14568));
    LocalMux I__1274 (
            .O(N__14568),
            .I(\PWMInstance7.un1_periodCounter12_1_0_a2_0_10 ));
    InMux I__1273 (
            .O(N__14565),
            .I(N__14562));
    LocalMux I__1272 (
            .O(N__14562),
            .I(\PWMInstance7.un1_periodCounter12_1_0_a2_0_9 ));
    CascadeMux I__1271 (
            .O(N__14559),
            .I(\PWMInstance7.un1_periodCounter12_1_0_a2_0_12_cascade_ ));
    InMux I__1270 (
            .O(N__14556),
            .I(N__14553));
    LocalMux I__1269 (
            .O(N__14553),
            .I(N__14550));
    Odrv4 I__1268 (
            .O(N__14550),
            .I(\PWMInstance7.un1_periodCounter12_1_0_a2_0_14 ));
    InMux I__1267 (
            .O(N__14547),
            .I(\PWMInstance7.un1_periodCounter_2_cry_10 ));
    InMux I__1266 (
            .O(N__14544),
            .I(\PWMInstance7.un1_periodCounter_2_cry_11 ));
    InMux I__1265 (
            .O(N__14541),
            .I(\PWMInstance7.un1_periodCounter_2_cry_12 ));
    InMux I__1264 (
            .O(N__14538),
            .I(\PWMInstance7.un1_periodCounter_2_cry_13 ));
    InMux I__1263 (
            .O(N__14535),
            .I(\PWMInstance7.un1_periodCounter_2_cry_14 ));
    InMux I__1262 (
            .O(N__14532),
            .I(bfn_2_10_0_));
    CascadeMux I__1261 (
            .O(N__14529),
            .I(N__14526));
    InMux I__1260 (
            .O(N__14526),
            .I(N__14521));
    InMux I__1259 (
            .O(N__14525),
            .I(N__14518));
    InMux I__1258 (
            .O(N__14524),
            .I(N__14515));
    LocalMux I__1257 (
            .O(N__14521),
            .I(N__14512));
    LocalMux I__1256 (
            .O(N__14518),
            .I(N__14509));
    LocalMux I__1255 (
            .O(N__14515),
            .I(\PWMInstance7.periodCounterZ0Z_16 ));
    Odrv4 I__1254 (
            .O(N__14512),
            .I(\PWMInstance7.periodCounterZ0Z_16 ));
    Odrv4 I__1253 (
            .O(N__14509),
            .I(\PWMInstance7.periodCounterZ0Z_16 ));
    CascadeMux I__1252 (
            .O(N__14502),
            .I(N__14498));
    InMux I__1251 (
            .O(N__14501),
            .I(N__14494));
    InMux I__1250 (
            .O(N__14498),
            .I(N__14491));
    InMux I__1249 (
            .O(N__14497),
            .I(N__14488));
    LocalMux I__1248 (
            .O(N__14494),
            .I(\PWMInstance7.periodCounter12 ));
    LocalMux I__1247 (
            .O(N__14491),
            .I(\PWMInstance7.periodCounter12 ));
    LocalMux I__1246 (
            .O(N__14488),
            .I(\PWMInstance7.periodCounter12 ));
    InMux I__1245 (
            .O(N__14481),
            .I(\PWMInstance7.un1_periodCounter_2_cry_1 ));
    InMux I__1244 (
            .O(N__14478),
            .I(\PWMInstance7.un1_periodCounter_2_cry_2 ));
    InMux I__1243 (
            .O(N__14475),
            .I(\PWMInstance7.un1_periodCounter_2_cry_3 ));
    InMux I__1242 (
            .O(N__14472),
            .I(\PWMInstance7.un1_periodCounter_2_cry_4 ));
    InMux I__1241 (
            .O(N__14469),
            .I(\PWMInstance7.un1_periodCounter_2_cry_5 ));
    InMux I__1240 (
            .O(N__14466),
            .I(\PWMInstance7.un1_periodCounter_2_cry_6 ));
    InMux I__1239 (
            .O(N__14463),
            .I(bfn_2_9_0_));
    InMux I__1238 (
            .O(N__14460),
            .I(\PWMInstance7.un1_periodCounter_2_cry_8 ));
    InMux I__1237 (
            .O(N__14457),
            .I(\PWMInstance7.un1_periodCounter_2_cry_9 ));
    IoInMux I__1236 (
            .O(N__14454),
            .I(N__14451));
    LocalMux I__1235 (
            .O(N__14451),
            .I(N__14448));
    IoSpan4Mux I__1234 (
            .O(N__14448),
            .I(N__14445));
    Odrv4 I__1233 (
            .O(N__14445),
            .I(CLK_c));
    CascadeMux I__1232 (
            .O(N__14442),
            .I(\PWMInstance7.un1_periodCounter12_1_0_a2_0_6_cascade_ ));
    InMux I__1231 (
            .O(N__14439),
            .I(\PWMInstance7.un1_periodCounter_2_cry_0 ));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(\QuadInstance7.un1_Quad_cry_7 ),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_12_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_5_0_));
    defparam IN_MUX_bfv_12_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_6_0_ (
            .carryinitin(\QuadInstance6.un1_Quad_cry_7 ),
            .carryinitout(bfn_12_6_0_));
    defparam IN_MUX_bfv_10_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_6_0_));
    defparam IN_MUX_bfv_10_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_7_0_ (
            .carryinitin(\QuadInstance5.un1_Quad_cry_7 ),
            .carryinitout(bfn_10_7_0_));
    defparam IN_MUX_bfv_15_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_3_0_));
    defparam IN_MUX_bfv_15_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_4_0_ (
            .carryinitin(\QuadInstance4.un1_Quad_cry_7 ),
            .carryinitout(bfn_15_4_0_));
    defparam IN_MUX_bfv_10_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_8_0_));
    defparam IN_MUX_bfv_10_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_9_0_ (
            .carryinitin(\QuadInstance3.un1_Quad_cry_7 ),
            .carryinitout(bfn_10_9_0_));
    defparam IN_MUX_bfv_7_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_6_0_));
    defparam IN_MUX_bfv_7_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_7_0_ (
            .carryinitin(\QuadInstance2.un1_Quad_cry_7 ),
            .carryinitout(bfn_7_7_0_));
    defparam IN_MUX_bfv_13_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_6_0_));
    defparam IN_MUX_bfv_13_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_7_0_ (
            .carryinitin(\QuadInstance1.un1_Quad_cry_7 ),
            .carryinitout(bfn_13_7_0_));
    defparam IN_MUX_bfv_17_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_6_0_));
    defparam IN_MUX_bfv_17_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_7_0_ (
            .carryinitin(\QuadInstance0.un1_Quad_cry_7 ),
            .carryinitout(bfn_17_7_0_));
    defparam IN_MUX_bfv_3_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_3_10_0_));
    defparam IN_MUX_bfv_3_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_3_11_0_ (
            .carryinitin(\PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_7 ),
            .carryinitout(bfn_3_11_0_));
    defparam IN_MUX_bfv_12_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_16_0_));
    defparam IN_MUX_bfv_12_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_17_0_ (
            .carryinitin(\PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_7 ),
            .carryinitout(bfn_12_17_0_));
    defparam IN_MUX_bfv_8_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_4_0_));
    defparam IN_MUX_bfv_8_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_5_0_ (
            .carryinitin(\PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_7 ),
            .carryinitout(bfn_8_5_0_));
    defparam IN_MUX_bfv_15_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_1_0_));
    defparam IN_MUX_bfv_15_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_2_0_ (
            .carryinitin(\PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_7 ),
            .carryinitout(bfn_15_2_0_));
    defparam IN_MUX_bfv_16_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_15_0_));
    defparam IN_MUX_bfv_16_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_16_0_ (
            .carryinitin(\PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_7 ),
            .carryinitout(bfn_16_16_0_));
    defparam IN_MUX_bfv_17_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_14_0_));
    defparam IN_MUX_bfv_17_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_15_0_ (
            .carryinitin(\PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_7 ),
            .carryinitout(bfn_17_15_0_));
    defparam IN_MUX_bfv_7_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_11_0_));
    defparam IN_MUX_bfv_7_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_12_0_ (
            .carryinitin(\PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_7 ),
            .carryinitout(bfn_7_12_0_));
    defparam IN_MUX_bfv_8_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_15_0_));
    defparam IN_MUX_bfv_8_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_16_0_ (
            .carryinitin(\PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_7 ),
            .carryinitout(bfn_8_16_0_));
    defparam IN_MUX_bfv_2_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_8_0_));
    defparam IN_MUX_bfv_2_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_9_0_ (
            .carryinitin(\PWMInstance7.un1_periodCounter_2_cry_7 ),
            .carryinitout(bfn_2_9_0_));
    defparam IN_MUX_bfv_2_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_10_0_ (
            .carryinitin(\PWMInstance7.un1_periodCounter_2_cry_15 ),
            .carryinitout(bfn_2_10_0_));
    defparam IN_MUX_bfv_11_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_14_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(\PWMInstance6.un1_periodCounter_2_cry_7 ),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_11_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_16_0_ (
            .carryinitin(\PWMInstance6.un1_periodCounter_2_cry_15 ),
            .carryinitout(bfn_11_16_0_));
    defparam IN_MUX_bfv_9_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_12_0_));
    defparam IN_MUX_bfv_9_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_13_0_ (
            .carryinitin(\PWMInstance5.un1_periodCounter_2_cry_7 ),
            .carryinitout(bfn_9_13_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(\PWMInstance5.un1_periodCounter_2_cry_15 ),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_14_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_16_0_));
    defparam IN_MUX_bfv_14_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_17_0_ (
            .carryinitin(\PWMInstance4.un1_periodCounter_2_cry_7 ),
            .carryinitout(bfn_14_17_0_));
    defparam IN_MUX_bfv_14_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_18_0_ (
            .carryinitin(\PWMInstance4.un1_periodCounter_2_cry_15 ),
            .carryinitout(bfn_14_18_0_));
    defparam IN_MUX_bfv_15_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_13_0_));
    defparam IN_MUX_bfv_15_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_14_0_ (
            .carryinitin(\PWMInstance3.un1_periodCounter_2_cry_7 ),
            .carryinitout(bfn_15_14_0_));
    defparam IN_MUX_bfv_15_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_15_0_ (
            .carryinitin(\PWMInstance3.un1_periodCounter_2_cry_15 ),
            .carryinitout(bfn_15_15_0_));
    defparam IN_MUX_bfv_18_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_11_0_));
    defparam IN_MUX_bfv_18_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_12_0_ (
            .carryinitin(\PWMInstance2.un1_periodCounter_2_cry_7 ),
            .carryinitout(bfn_18_12_0_));
    defparam IN_MUX_bfv_18_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_13_0_ (
            .carryinitin(\PWMInstance2.un1_periodCounter_2_cry_15 ),
            .carryinitout(bfn_18_13_0_));
    defparam IN_MUX_bfv_8_1_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_1_0_));
    defparam IN_MUX_bfv_8_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_2_0_ (
            .carryinitin(\PWMInstance1.un1_periodCounter_2_cry_7 ),
            .carryinitout(bfn_8_2_0_));
    defparam IN_MUX_bfv_8_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_3_0_ (
            .carryinitin(\PWMInstance1.un1_periodCounter_2_cry_15 ),
            .carryinitout(bfn_8_3_0_));
    defparam IN_MUX_bfv_7_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_16_0_));
    defparam IN_MUX_bfv_7_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_17_0_ (
            .carryinitin(\PWMInstance0.un1_periodCounter_2_cry_7 ),
            .carryinitout(bfn_7_17_0_));
    defparam IN_MUX_bfv_7_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_18_0_ (
            .carryinitin(\PWMInstance0.un1_periodCounter_2_cry_15 ),
            .carryinitout(bfn_7_18_0_));
    SMCCLK internalOscilator (
            .CLK(internalOscilatorOutputNet));
    ICE_GB SCKr_RNIBA7C_0_2 (
            .USERSIGNALTOGLOBALBUFFER(N__37941),
            .GLOBALBUFFEROUTPUT(N_1187_g));
    ICE_GB SCKr_RNIMKEO_0_2 (
            .USERSIGNALTOGLOBALBUFFER(N__37923),
            .GLOBALBUFFEROUTPUT(N_45_0_g));
    ICE_GB RST_ibuf_RNIUR47_0 (
            .USERSIGNALTOGLOBALBUFFER(N__15207),
            .GLOBALBUFFEROUTPUT(RST_c_i_g));
    ICE_GB \PWMInstance0.N_42_g_gb  (
            .USERSIGNALTOGLOBALBUFFER(N__25626),
            .GLOBALBUFFEROUTPUT(PWMInstance0_N_42_g));
    ICE_GB My_Global_Buffer_i (
            .USERSIGNALTOGLOBALBUFFER(N__14454),
            .GLOBALBUFFEROUTPUT(myclk));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \PWMInstance7.periodCounter_RNIG0CG_16_LC_2_7_6 .C_ON=1'b0;
    defparam \PWMInstance7.periodCounter_RNIG0CG_16_LC_2_7_6 .SEQ_MODE=4'b0000;
    defparam \PWMInstance7.periodCounter_RNIG0CG_16_LC_2_7_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \PWMInstance7.periodCounter_RNIG0CG_16_LC_2_7_6  (
            .in0(_gnd_net_),
            .in1(N__14525),
            .in2(_gnd_net_),
            .in3(N__14971),
            .lcout(),
            .ltout(\PWMInstance7.un1_periodCounter12_1_0_a2_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance7.periodCounter_RNI7VP12_1_LC_2_7_7 .C_ON=1'b0;
    defparam \PWMInstance7.periodCounter_RNI7VP12_1_LC_2_7_7 .SEQ_MODE=4'b0000;
    defparam \PWMInstance7.periodCounter_RNI7VP12_1_LC_2_7_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \PWMInstance7.periodCounter_RNI7VP12_1_LC_2_7_7  (
            .in0(N__14842),
            .in1(N__15028),
            .in2(N__14442),
            .in3(N__14497),
            .lcout(\PWMInstance7.un1_periodCounter12_1_0_a2_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance7.periodCounter_0_LC_2_8_0 .C_ON=1'b1;
    defparam \PWMInstance7.periodCounter_0_LC_2_8_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.periodCounter_0_LC_2_8_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance7.periodCounter_0_LC_2_8_0  (
            .in0(_gnd_net_),
            .in1(N__15055),
            .in2(N__14502),
            .in3(N__14501),
            .lcout(\PWMInstance7.periodCounterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_2_8_0_),
            .carryout(\PWMInstance7.un1_periodCounter_2_cry_0 ),
            .clk(N__38625),
            .ce(),
            .sr(N__35314));
    defparam \PWMInstance7.periodCounter_1_LC_2_8_1 .C_ON=1'b1;
    defparam \PWMInstance7.periodCounter_1_LC_2_8_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.periodCounter_1_LC_2_8_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance7.periodCounter_1_LC_2_8_1  (
            .in0(_gnd_net_),
            .in1(N__15029),
            .in2(_gnd_net_),
            .in3(N__14439),
            .lcout(\PWMInstance7.periodCounterZ0Z_1 ),
            .ltout(),
            .carryin(\PWMInstance7.un1_periodCounter_2_cry_0 ),
            .carryout(\PWMInstance7.un1_periodCounter_2_cry_1 ),
            .clk(N__38625),
            .ce(),
            .sr(N__35314));
    defparam \PWMInstance7.periodCounter_2_LC_2_8_2 .C_ON=1'b1;
    defparam \PWMInstance7.periodCounter_2_LC_2_8_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.periodCounter_2_LC_2_8_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance7.periodCounter_2_LC_2_8_2  (
            .in0(_gnd_net_),
            .in1(N__14652),
            .in2(_gnd_net_),
            .in3(N__14481),
            .lcout(\PWMInstance7.periodCounterZ0Z_2 ),
            .ltout(),
            .carryin(\PWMInstance7.un1_periodCounter_2_cry_1 ),
            .carryout(\PWMInstance7.un1_periodCounter_2_cry_2 ),
            .clk(N__38625),
            .ce(),
            .sr(N__35314));
    defparam \PWMInstance7.periodCounter_3_LC_2_8_3 .C_ON=1'b1;
    defparam \PWMInstance7.periodCounter_3_LC_2_8_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.periodCounter_3_LC_2_8_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance7.periodCounter_3_LC_2_8_3  (
            .in0(_gnd_net_),
            .in1(N__14636),
            .in2(_gnd_net_),
            .in3(N__14478),
            .lcout(\PWMInstance7.periodCounterZ0Z_3 ),
            .ltout(),
            .carryin(\PWMInstance7.un1_periodCounter_2_cry_2 ),
            .carryout(\PWMInstance7.un1_periodCounter_2_cry_3 ),
            .clk(N__38625),
            .ce(),
            .sr(N__35314));
    defparam \PWMInstance7.periodCounter_4_LC_2_8_4 .C_ON=1'b1;
    defparam \PWMInstance7.periodCounter_4_LC_2_8_4 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.periodCounter_4_LC_2_8_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance7.periodCounter_4_LC_2_8_4  (
            .in0(_gnd_net_),
            .in1(N__14787),
            .in2(_gnd_net_),
            .in3(N__14475),
            .lcout(\PWMInstance7.periodCounterZ0Z_4 ),
            .ltout(),
            .carryin(\PWMInstance7.un1_periodCounter_2_cry_3 ),
            .carryout(\PWMInstance7.un1_periodCounter_2_cry_4 ),
            .clk(N__38625),
            .ce(),
            .sr(N__35314));
    defparam \PWMInstance7.periodCounter_5_LC_2_8_5 .C_ON=1'b1;
    defparam \PWMInstance7.periodCounter_5_LC_2_8_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.periodCounter_5_LC_2_8_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance7.periodCounter_5_LC_2_8_5  (
            .in0(_gnd_net_),
            .in1(N__14771),
            .in2(_gnd_net_),
            .in3(N__14472),
            .lcout(\PWMInstance7.periodCounterZ0Z_5 ),
            .ltout(),
            .carryin(\PWMInstance7.un1_periodCounter_2_cry_4 ),
            .carryout(\PWMInstance7.un1_periodCounter_2_cry_5 ),
            .clk(N__38625),
            .ce(),
            .sr(N__35314));
    defparam \PWMInstance7.periodCounter_6_LC_2_8_6 .C_ON=1'b1;
    defparam \PWMInstance7.periodCounter_6_LC_2_8_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.periodCounter_6_LC_2_8_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance7.periodCounter_6_LC_2_8_6  (
            .in0(_gnd_net_),
            .in1(N__14999),
            .in2(_gnd_net_),
            .in3(N__14469),
            .lcout(\PWMInstance7.periodCounterZ0Z_6 ),
            .ltout(),
            .carryin(\PWMInstance7.un1_periodCounter_2_cry_5 ),
            .carryout(\PWMInstance7.un1_periodCounter_2_cry_6 ),
            .clk(N__38625),
            .ce(),
            .sr(N__35314));
    defparam \PWMInstance7.periodCounter_7_LC_2_8_7 .C_ON=1'b1;
    defparam \PWMInstance7.periodCounter_7_LC_2_8_7 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.periodCounter_7_LC_2_8_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance7.periodCounter_7_LC_2_8_7  (
            .in0(N__14929),
            .in1(N__14975),
            .in2(_gnd_net_),
            .in3(N__14466),
            .lcout(\PWMInstance7.periodCounterZ0Z_7 ),
            .ltout(),
            .carryin(\PWMInstance7.un1_periodCounter_2_cry_6 ),
            .carryout(\PWMInstance7.un1_periodCounter_2_cry_7 ),
            .clk(N__38625),
            .ce(),
            .sr(N__35314));
    defparam \PWMInstance7.periodCounter_8_LC_2_9_0 .C_ON=1'b1;
    defparam \PWMInstance7.periodCounter_8_LC_2_9_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.periodCounter_8_LC_2_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance7.periodCounter_8_LC_2_9_0  (
            .in0(_gnd_net_),
            .in1(N__14754),
            .in2(_gnd_net_),
            .in3(N__14463),
            .lcout(\PWMInstance7.periodCounterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_2_9_0_),
            .carryout(\PWMInstance7.un1_periodCounter_2_cry_8 ),
            .clk(N__38614),
            .ce(),
            .sr(N__35312));
    defparam \PWMInstance7.periodCounter_9_LC_2_9_1 .C_ON=1'b1;
    defparam \PWMInstance7.periodCounter_9_LC_2_9_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.periodCounter_9_LC_2_9_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance7.periodCounter_9_LC_2_9_1  (
            .in0(_gnd_net_),
            .in1(N__14738),
            .in2(_gnd_net_),
            .in3(N__14460),
            .lcout(\PWMInstance7.periodCounterZ0Z_9 ),
            .ltout(),
            .carryin(\PWMInstance7.un1_periodCounter_2_cry_8 ),
            .carryout(\PWMInstance7.un1_periodCounter_2_cry_9 ),
            .clk(N__38614),
            .ce(),
            .sr(N__35312));
    defparam \PWMInstance7.periodCounter_10_LC_2_9_2 .C_ON=1'b1;
    defparam \PWMInstance7.periodCounter_10_LC_2_9_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.periodCounter_10_LC_2_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance7.periodCounter_10_LC_2_9_2  (
            .in0(_gnd_net_),
            .in1(N__14596),
            .in2(_gnd_net_),
            .in3(N__14457),
            .lcout(\PWMInstance7.periodCounterZ0Z_10 ),
            .ltout(),
            .carryin(\PWMInstance7.un1_periodCounter_2_cry_9 ),
            .carryout(\PWMInstance7.un1_periodCounter_2_cry_10 ),
            .clk(N__38614),
            .ce(),
            .sr(N__35312));
    defparam \PWMInstance7.periodCounter_11_LC_2_9_3 .C_ON=1'b1;
    defparam \PWMInstance7.periodCounter_11_LC_2_9_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.periodCounter_11_LC_2_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance7.periodCounter_11_LC_2_9_3  (
            .in0(N__14938),
            .in1(N__14615),
            .in2(_gnd_net_),
            .in3(N__14547),
            .lcout(\PWMInstance7.periodCounterZ0Z_11 ),
            .ltout(),
            .carryin(\PWMInstance7.un1_periodCounter_2_cry_10 ),
            .carryout(\PWMInstance7.un1_periodCounter_2_cry_11 ),
            .clk(N__38614),
            .ce(),
            .sr(N__35312));
    defparam \PWMInstance7.periodCounter_12_LC_2_9_4 .C_ON=1'b1;
    defparam \PWMInstance7.periodCounter_12_LC_2_9_4 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.periodCounter_12_LC_2_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance7.periodCounter_12_LC_2_9_4  (
            .in0(N__14927),
            .in1(N__15118),
            .in2(_gnd_net_),
            .in3(N__14544),
            .lcout(\PWMInstance7.periodCounterZ0Z_12 ),
            .ltout(),
            .carryin(\PWMInstance7.un1_periodCounter_2_cry_11 ),
            .carryout(\PWMInstance7.un1_periodCounter_2_cry_12 ),
            .clk(N__38614),
            .ce(),
            .sr(N__35312));
    defparam \PWMInstance7.periodCounter_13_LC_2_9_5 .C_ON=1'b1;
    defparam \PWMInstance7.periodCounter_13_LC_2_9_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.periodCounter_13_LC_2_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance7.periodCounter_13_LC_2_9_5  (
            .in0(N__14939),
            .in1(N__15088),
            .in2(_gnd_net_),
            .in3(N__14541),
            .lcout(\PWMInstance7.periodCounterZ0Z_13 ),
            .ltout(),
            .carryin(\PWMInstance7.un1_periodCounter_2_cry_12 ),
            .carryout(\PWMInstance7.un1_periodCounter_2_cry_13 ),
            .clk(N__38614),
            .ce(),
            .sr(N__35312));
    defparam \PWMInstance7.periodCounter_14_LC_2_9_6 .C_ON=1'b1;
    defparam \PWMInstance7.periodCounter_14_LC_2_9_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.periodCounter_14_LC_2_9_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance7.periodCounter_14_LC_2_9_6  (
            .in0(_gnd_net_),
            .in1(N__14820),
            .in2(_gnd_net_),
            .in3(N__14538),
            .lcout(\PWMInstance7.periodCounterZ0Z_14 ),
            .ltout(),
            .carryin(\PWMInstance7.un1_periodCounter_2_cry_13 ),
            .carryout(\PWMInstance7.un1_periodCounter_2_cry_14 ),
            .clk(N__38614),
            .ce(),
            .sr(N__35312));
    defparam \PWMInstance7.periodCounter_15_LC_2_9_7 .C_ON=1'b1;
    defparam \PWMInstance7.periodCounter_15_LC_2_9_7 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.periodCounter_15_LC_2_9_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance7.periodCounter_15_LC_2_9_7  (
            .in0(_gnd_net_),
            .in1(N__14844),
            .in2(_gnd_net_),
            .in3(N__14535),
            .lcout(\PWMInstance7.periodCounterZ0Z_15 ),
            .ltout(),
            .carryin(\PWMInstance7.un1_periodCounter_2_cry_14 ),
            .carryout(\PWMInstance7.un1_periodCounter_2_cry_15 ),
            .clk(N__38614),
            .ce(),
            .sr(N__35312));
    defparam \PWMInstance7.periodCounter_16_LC_2_10_0 .C_ON=1'b0;
    defparam \PWMInstance7.periodCounter_16_LC_2_10_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.periodCounter_16_LC_2_10_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance7.periodCounter_16_LC_2_10_0  (
            .in0(N__14928),
            .in1(N__14524),
            .in2(_gnd_net_),
            .in3(N__14532),
            .lcout(\PWMInstance7.periodCounterZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38603),
            .ce(),
            .sr(N__35311));
    defparam \PWMInstance7.out_RNO_0_LC_3_7_0 .C_ON=1'b0;
    defparam \PWMInstance7.out_RNO_0_LC_3_7_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance7.out_RNO_0_LC_3_7_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \PWMInstance7.out_RNO_0_LC_3_7_0  (
            .in0(N__14871),
            .in1(N__14671),
            .in2(N__14529),
            .in3(N__14692),
            .lcout(\PWMInstance7.un1_periodCounter12_1_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance7.clkCount_0_LC_3_7_1 .C_ON=1'b0;
    defparam \PWMInstance7.clkCount_0_LC_3_7_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.clkCount_0_LC_3_7_1 .LUT_INIT=16'b1010101000000101;
    LogicCell40 \PWMInstance7.clkCount_0_LC_3_7_1  (
            .in0(N__14693),
            .in1(_gnd_net_),
            .in2(N__14678),
            .in3(N__17813),
            .lcout(\PWMInstance7.clkCountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38626),
            .ce(),
            .sr(N__35695));
    defparam \PWMInstance7.clkCount_RNIE5211_0_LC_3_7_2 .C_ON=1'b0;
    defparam \PWMInstance7.clkCount_RNIE5211_0_LC_3_7_2 .SEQ_MODE=4'b0000;
    defparam \PWMInstance7.clkCount_RNIE5211_0_LC_3_7_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \PWMInstance7.clkCount_RNIE5211_0_LC_3_7_2  (
            .in0(N__14870),
            .in1(N__14670),
            .in2(_gnd_net_),
            .in3(N__14691),
            .lcout(\PWMInstance7.periodCounter12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance7.clkCount_1_LC_3_7_3 .C_ON=1'b0;
    defparam \PWMInstance7.clkCount_1_LC_3_7_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.clkCount_1_LC_3_7_3 .LUT_INIT=16'b1111000000001010;
    LogicCell40 \PWMInstance7.clkCount_1_LC_3_7_3  (
            .in0(N__14694),
            .in1(_gnd_net_),
            .in2(N__14679),
            .in3(N__17814),
            .lcout(\PWMInstance7.clkCountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38626),
            .ce(),
            .sr(N__35695));
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_3_8_1 .C_ON=1'b0;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_3_8_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_3_8_1 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \PWMInstance7.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_3_8_1  (
            .in0(N__14651),
            .in1(N__14850),
            .in2(N__14637),
            .in3(N__14658),
            .lcout(\PWMInstance7.un1_PWMPulseWidthCount_0_I_9_c_RNO_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance7.PWMPulseWidthCount_esr_2_LC_3_8_2 .C_ON=1'b0;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_2_LC_3_8_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_2_LC_3_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance7.PWMPulseWidthCount_esr_2_LC_3_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31604),
            .lcout(\PWMInstance7.PWMPulseWidthCountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38615),
            .ce(N__15270),
            .sr(N__35702));
    defparam \PWMInstance7.periodCounter_RNI9PBG_2_LC_3_8_4 .C_ON=1'b0;
    defparam \PWMInstance7.periodCounter_RNI9PBG_2_LC_3_8_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance7.periodCounter_RNI9PBG_2_LC_3_8_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \PWMInstance7.periodCounter_RNI9PBG_2_LC_3_8_4  (
            .in0(_gnd_net_),
            .in1(N__14812),
            .in2(_gnd_net_),
            .in3(N__14650),
            .lcout(\PWMInstance7.un1_periodCounter12_1_0_a2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance7.periodCounter_RNI79MR_3_LC_3_9_0 .C_ON=1'b0;
    defparam \PWMInstance7.periodCounter_RNI79MR_3_LC_3_9_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance7.periodCounter_RNI79MR_3_LC_3_9_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \PWMInstance7.periodCounter_RNI79MR_3_LC_3_9_0  (
            .in0(N__14737),
            .in1(N__14770),
            .in2(N__14616),
            .in3(N__14635),
            .lcout(\PWMInstance7.un1_periodCounter12_1_0_a2_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_3_9_1 .C_ON=1'b0;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_3_9_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_3_9_1 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \PWMInstance7.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_3_9_1  (
            .in0(N__15180),
            .in1(N__14611),
            .in2(N__14597),
            .in3(N__14856),
            .lcout(\PWMInstance7.un1_PWMPulseWidthCount_0_I_33_c_RNO_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance7.periodCounter_RNI68MR_0_LC_3_9_2 .C_ON=1'b0;
    defparam \PWMInstance7.periodCounter_RNI68MR_0_LC_3_9_2 .SEQ_MODE=4'b0000;
    defparam \PWMInstance7.periodCounter_RNI68MR_0_LC_3_9_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \PWMInstance7.periodCounter_RNI68MR_0_LC_3_9_2  (
            .in0(N__14753),
            .in1(N__14998),
            .in2(N__15095),
            .in3(N__15056),
            .lcout(\PWMInstance7.un1_periodCounter12_1_0_a2_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance7.periodCounter_RNIS3EB1_4_LC_3_9_3 .C_ON=1'b0;
    defparam \PWMInstance7.periodCounter_RNIS3EB1_4_LC_3_9_3 .SEQ_MODE=4'b0000;
    defparam \PWMInstance7.periodCounter_RNIS3EB1_4_LC_3_9_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \PWMInstance7.periodCounter_RNIS3EB1_4_LC_3_9_3  (
            .in0(N__14786),
            .in1(N__15120),
            .in2(N__14598),
            .in3(N__14577),
            .lcout(),
            .ltout(\PWMInstance7.un1_periodCounter12_1_0_a2_0_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance7.periodCounter_RNIGKK45_0_LC_3_9_4 .C_ON=1'b0;
    defparam \PWMInstance7.periodCounter_RNIGKK45_0_LC_3_9_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance7.periodCounter_RNIGKK45_0_LC_3_9_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \PWMInstance7.periodCounter_RNIGKK45_0_LC_3_9_4  (
            .in0(N__14571),
            .in1(N__14565),
            .in2(N__14559),
            .in3(N__14556),
            .lcout(\PWMInstance7.out_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_3_9_5 .C_ON=1'b0;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_3_9_5 .SEQ_MODE=4'b0000;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_3_9_5 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \PWMInstance7.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_3_9_5  (
            .in0(N__14785),
            .in1(N__15165),
            .in2(N__14772),
            .in3(N__15156),
            .lcout(\PWMInstance7.un1_PWMPulseWidthCount_0_I_15_c_RNO_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_3_9_6 .C_ON=1'b0;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_3_9_6 .SEQ_MODE=4'b0000;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_3_9_6 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \PWMInstance7.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_3_9_6  (
            .in0(N__14752),
            .in1(N__14862),
            .in2(N__14739),
            .in3(N__15195),
            .lcout(\PWMInstance7.un1_PWMPulseWidthCount_0_I_45_c_RNO_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_1_c_LC_3_10_0 .C_ON=1'b1;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_1_c_LC_3_10_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_1_c_LC_3_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance7.un1_PWMPulseWidthCount_0_I_1_c_LC_3_10_0  (
            .in0(_gnd_net_),
            .in1(N__15009),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_3_10_0_),
            .carryout(\PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_9_c_LC_3_10_1 .C_ON=1'b1;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_9_c_LC_3_10_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_9_c_LC_3_10_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance7.un1_PWMPulseWidthCount_0_I_9_c_LC_3_10_1  (
            .in0(_gnd_net_),
            .in1(N__14721),
            .in2(N__32585),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_0 ),
            .carryout(\PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_15_c_LC_3_10_2 .C_ON=1'b1;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_15_c_LC_3_10_2 .SEQ_MODE=4'b0000;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_15_c_LC_3_10_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance7.un1_PWMPulseWidthCount_0_I_15_c_LC_3_10_2  (
            .in0(_gnd_net_),
            .in1(N__14712),
            .in2(N__32580),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_1 ),
            .carryout(\PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_27_c_LC_3_10_3 .C_ON=1'b1;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_27_c_LC_3_10_3 .SEQ_MODE=4'b0000;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_27_c_LC_3_10_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance7.un1_PWMPulseWidthCount_0_I_27_c_LC_3_10_3  (
            .in0(_gnd_net_),
            .in1(N__14955),
            .in2(N__32583),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_2 ),
            .carryout(\PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_45_c_LC_3_10_4 .C_ON=1'b1;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_45_c_LC_3_10_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_45_c_LC_3_10_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance7.un1_PWMPulseWidthCount_0_I_45_c_LC_3_10_4  (
            .in0(_gnd_net_),
            .in1(N__14706),
            .in2(N__32581),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_3 ),
            .carryout(\PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_33_c_LC_3_10_5 .C_ON=1'b1;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_33_c_LC_3_10_5 .SEQ_MODE=4'b0000;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_33_c_LC_3_10_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance7.un1_PWMPulseWidthCount_0_I_33_c_LC_3_10_5  (
            .in0(_gnd_net_),
            .in1(N__14700),
            .in2(N__32584),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_4 ),
            .carryout(\PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_39_c_LC_3_10_6 .C_ON=1'b1;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_39_c_LC_3_10_6 .SEQ_MODE=4'b0000;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_39_c_LC_3_10_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance7.un1_PWMPulseWidthCount_0_I_39_c_LC_3_10_6  (
            .in0(_gnd_net_),
            .in1(N__32534),
            .in2(N__15069),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_5 ),
            .carryout(\PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_21_c_LC_3_10_7 .C_ON=1'b1;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_21_c_LC_3_10_7 .SEQ_MODE=4'b0000;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_21_c_LC_3_10_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance7.un1_PWMPulseWidthCount_0_I_21_c_LC_3_10_7  (
            .in0(_gnd_net_),
            .in1(N__14799),
            .in2(N__32582),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_6 ),
            .carryout(\PWMInstance7.un1_PWMPulseWidthCount_0_data_tmp_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance7.out_LC_3_11_0 .C_ON=1'b0;
    defparam \PWMInstance7.out_LC_3_11_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.out_LC_3_11_0 .LUT_INIT=16'b1111101011110010;
    LogicCell40 \PWMInstance7.out_LC_3_11_0  (
            .in0(N__14882),
            .in1(N__14949),
            .in2(N__14940),
            .in3(N__14898),
            .lcout(PWM7_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38585),
            .ce(),
            .sr(N__35726));
    defparam pwmWrite_fast_7_LC_4_7_0.C_ON=1'b0;
    defparam pwmWrite_fast_7_LC_4_7_0.SEQ_MODE=4'b1000;
    defparam pwmWrite_fast_7_LC_4_7_0.LUT_INIT=16'b0000100000000000;
    LogicCell40 pwmWrite_fast_7_LC_4_7_0 (
            .in0(N__33857),
            .in1(N__33670),
            .in2(N__33449),
            .in3(N__23463),
            .lcout(pwmWrite_fastZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38616),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance7.PWMPulseWidthCount_esr_9_LC_4_8_3 .C_ON=1'b0;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_9_LC_4_8_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_9_LC_4_8_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \PWMInstance7.PWMPulseWidthCount_esr_9_LC_4_8_3  (
            .in0(N__28580),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PWMInstance7.PWMPulseWidthCountZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38604),
            .ce(N__15266),
            .sr(N__35696));
    defparam \PWMInstance7.PWMPulseWidthCount_esr_10_LC_4_8_5 .C_ON=1'b0;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_10_LC_4_8_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_10_LC_4_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance7.PWMPulseWidthCount_esr_10_LC_4_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36167),
            .lcout(\PWMInstance7.PWMPulseWidthCountZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38604),
            .ce(N__15266),
            .sr(N__35696));
    defparam \PWMInstance7.PWMPulseWidthCount_esr_3_LC_4_8_7 .C_ON=1'b0;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_3_LC_4_8_7 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_3_LC_4_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance7.PWMPulseWidthCount_esr_3_LC_4_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32084),
            .lcout(\PWMInstance7.PWMPulseWidthCountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38604),
            .ce(N__15266),
            .sr(N__35696));
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_4_9_0 .C_ON=1'b0;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_4_9_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \PWMInstance7.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_4_9_0  (
            .in0(N__14793),
            .in1(N__14843),
            .in2(N__15129),
            .in3(N__14819),
            .lcout(\PWMInstance7.un1_PWMPulseWidthCount_0_I_21_c_RNO_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance7.PWMPulseWidthCount_esr_14_LC_4_9_1 .C_ON=1'b0;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_14_LC_4_9_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_14_LC_4_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance7.PWMPulseWidthCount_esr_14_LC_4_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34399),
            .lcout(\PWMInstance7.PWMPulseWidthCountZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38595),
            .ce(N__15279),
            .sr(N__35703));
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_4_9_6 .C_ON=1'b0;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_4_9_6 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \PWMInstance7.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_4_9_6  (
            .in0(N__15171),
            .in1(N__15119),
            .in2(N__15096),
            .in3(N__15186),
            .lcout(\PWMInstance7.un1_PWMPulseWidthCount_0_I_39_c_RNO_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_4_10_1 .C_ON=1'b0;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_4_10_1 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance7.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_4_10_1  (
            .in0(N__15294),
            .in1(N__15060),
            .in2(N__15036),
            .in3(N__15285),
            .lcout(\PWMInstance7.un1_PWMPulseWidthCount_0_I_1_c_RNO_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_4_10_4 .C_ON=1'b0;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance7.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_4_10_4 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \PWMInstance7.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_4_10_4  (
            .in0(N__15003),
            .in1(N__15138),
            .in2(N__15147),
            .in3(N__14979),
            .lcout(\PWMInstance7.un1_PWMPulseWidthCount_0_I_27_c_RNO_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.PWMPulseWidthCount_esr_10_LC_4_13_3 .C_ON=1'b0;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_10_LC_4_13_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_10_LC_4_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance5.PWMPulseWidthCount_esr_10_LC_4_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36166),
            .lcout(\PWMInstance5.PWMPulseWidthCountZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38557),
            .ce(N__19651),
            .sr(N__35736));
    defparam \PWMInstance5.PWMPulseWidthCount_esr_9_LC_4_14_6 .C_ON=1'b0;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_9_LC_4_14_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_9_LC_4_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance5.PWMPulseWidthCount_esr_9_LC_4_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28579),
            .lcout(\PWMInstance5.PWMPulseWidthCountZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38551),
            .ce(N__19653),
            .sr(N__35741));
    defparam \PWMInstance1.PWMPulseWidthCount_esr_8_LC_5_4_0 .C_ON=1'b0;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_8_LC_5_4_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_8_LC_5_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance1.PWMPulseWidthCount_esr_8_LC_5_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29007),
            .lcout(\PWMInstance1.PWMPulseWidthCountZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38637),
            .ce(N__16826),
            .sr(N__35678));
    defparam \PWMInstance1.PWMPulseWidthCount_esr_7_LC_5_4_1 .C_ON=1'b0;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_7_LC_5_4_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_7_LC_5_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance1.PWMPulseWidthCount_esr_7_LC_5_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29417),
            .lcout(\PWMInstance1.PWMPulseWidthCountZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38637),
            .ce(N__16826),
            .sr(N__35678));
    defparam \PWMInstance1.PWMPulseWidthCount_esr_11_LC_5_4_3 .C_ON=1'b0;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_11_LC_5_4_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_11_LC_5_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance1.PWMPulseWidthCount_esr_11_LC_5_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36003),
            .lcout(\PWMInstance1.PWMPulseWidthCountZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38637),
            .ce(N__16826),
            .sr(N__35678));
    defparam \PWMInstance1.PWMPulseWidthCount_esr_14_LC_5_7_7 .C_ON=1'b0;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_14_LC_5_7_7 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_14_LC_5_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance1.PWMPulseWidthCount_esr_14_LC_5_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34414),
            .lcout(\PWMInstance1.PWMPulseWidthCountZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38605),
            .ce(N__16822),
            .sr(N__35683));
    defparam \PWMInstance7.PWMPulseWidthCount_esr_ctle_15_LC_5_8_4 .C_ON=1'b0;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_ctle_15_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_ctle_15_LC_5_8_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \PWMInstance7.PWMPulseWidthCount_esr_ctle_15_LC_5_8_4  (
            .in0(N__35824),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17807),
            .lcout(\PWMInstance7.pwmWrite_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance7.PWMPulseWidthCount_esr_8_LC_5_9_0 .C_ON=1'b0;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_8_LC_5_9_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_8_LC_5_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance7.PWMPulseWidthCount_esr_8_LC_5_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29003),
            .lcout(\PWMInstance7.PWMPulseWidthCountZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38586),
            .ce(N__15275),
            .sr(N__35697));
    defparam \PWMInstance7.PWMPulseWidthCount_esr_13_LC_5_9_2 .C_ON=1'b0;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_13_LC_5_9_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_13_LC_5_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance7.PWMPulseWidthCount_esr_13_LC_5_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28725),
            .lcout(\PWMInstance7.PWMPulseWidthCountZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38586),
            .ce(N__15275),
            .sr(N__35697));
    defparam \PWMInstance7.PWMPulseWidthCount_esr_11_LC_5_9_3 .C_ON=1'b0;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_11_LC_5_9_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_11_LC_5_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance7.PWMPulseWidthCount_esr_11_LC_5_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36002),
            .lcout(\PWMInstance7.PWMPulseWidthCountZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38586),
            .ce(N__15275),
            .sr(N__35697));
    defparam \PWMInstance7.PWMPulseWidthCount_esr_12_LC_5_9_4 .C_ON=1'b0;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_12_LC_5_9_4 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_12_LC_5_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance7.PWMPulseWidthCount_esr_12_LC_5_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28873),
            .lcout(\PWMInstance7.PWMPulseWidthCountZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38586),
            .ce(N__15275),
            .sr(N__35697));
    defparam \PWMInstance7.PWMPulseWidthCount_esr_5_LC_5_9_5 .C_ON=1'b0;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_5_LC_5_9_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_5_LC_5_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance7.PWMPulseWidthCount_esr_5_LC_5_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36376),
            .lcout(\PWMInstance7.PWMPulseWidthCountZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38586),
            .ce(N__15275),
            .sr(N__35697));
    defparam \PWMInstance7.PWMPulseWidthCount_esr_4_LC_5_9_7 .C_ON=1'b0;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_4_LC_5_9_7 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_4_LC_5_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance7.PWMPulseWidthCount_esr_4_LC_5_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36503),
            .lcout(\PWMInstance7.PWMPulseWidthCountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38586),
            .ce(N__15275),
            .sr(N__35697));
    defparam \PWMInstance7.PWMPulseWidthCount_esr_7_LC_5_10_0 .C_ON=1'b0;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_7_LC_5_10_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_7_LC_5_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance7.PWMPulseWidthCount_esr_7_LC_5_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29460),
            .lcout(\PWMInstance7.PWMPulseWidthCountZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38574),
            .ce(N__15271),
            .sr(N__35704));
    defparam \PWMInstance7.PWMPulseWidthCount_esr_6_LC_5_10_2 .C_ON=1'b0;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_6_LC_5_10_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_6_LC_5_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance7.PWMPulseWidthCount_esr_6_LC_5_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31125),
            .lcout(\PWMInstance7.PWMPulseWidthCountZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38574),
            .ce(N__15271),
            .sr(N__35704));
    defparam \PWMInstance7.PWMPulseWidthCount_esr_15_LC_5_10_5 .C_ON=1'b0;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_15_LC_5_10_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_15_LC_5_10_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \PWMInstance7.PWMPulseWidthCount_esr_15_LC_5_10_5  (
            .in0(N__31894),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PWMInstance7.PWMPulseWidthCountZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38574),
            .ce(N__15271),
            .sr(N__35704));
    defparam \PWMInstance7.PWMPulseWidthCount_esr_1_LC_5_10_6 .C_ON=1'b0;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_1_LC_5_10_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_1_LC_5_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance7.PWMPulseWidthCount_esr_1_LC_5_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31278),
            .lcout(\PWMInstance7.PWMPulseWidthCountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38574),
            .ce(N__15271),
            .sr(N__35704));
    defparam \PWMInstance7.PWMPulseWidthCount_esr_0_LC_5_10_7 .C_ON=1'b0;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_0_LC_5_10_7 .SEQ_MODE=4'b1000;
    defparam \PWMInstance7.PWMPulseWidthCount_esr_0_LC_5_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance7.PWMPulseWidthCount_esr_0_LC_5_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31436),
            .lcout(\PWMInstance7.PWMPulseWidthCountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38574),
            .ce(N__15271),
            .sr(N__35704));
    defparam \PWMInstance0.PWMPulseWidthCount_esr_10_LC_5_11_3 .C_ON=1'b0;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_10_LC_5_11_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_10_LC_5_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance0.PWMPulseWidthCount_esr_10_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36149),
            .lcout(\PWMInstance0.PWMPulseWidthCountZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38565),
            .ce(N__18249),
            .sr(N__35708));
    defparam \PWMInstance5.PWMPulseWidthCount_esr_8_LC_5_12_2 .C_ON=1'b0;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_8_LC_5_12_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_8_LC_5_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance5.PWMPulseWidthCount_esr_8_LC_5_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29002),
            .lcout(\PWMInstance5.PWMPulseWidthCountZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38558),
            .ce(N__19650),
            .sr(N__35718));
    defparam \PWMInstance5.PWMPulseWidthCount_esr_14_LC_5_12_3 .C_ON=1'b0;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_14_LC_5_12_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_14_LC_5_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance5.PWMPulseWidthCount_esr_14_LC_5_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34413),
            .lcout(\PWMInstance5.PWMPulseWidthCountZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38558),
            .ce(N__19650),
            .sr(N__35718));
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_5_13_3 .C_ON=1'b0;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_5_13_3 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \PWMInstance5.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_5_13_3  (
            .in0(N__17942),
            .in1(N__15219),
            .in2(N__19419),
            .in3(N__15213),
            .lcout(\PWMInstance5.un1_PWMPulseWidthCount_0_I_45_c_RNO_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.PWMPulseWidthCount_esr_12_LC_5_14_2 .C_ON=1'b0;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_12_LC_5_14_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_12_LC_5_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance5.PWMPulseWidthCount_esr_12_LC_5_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28872),
            .lcout(\PWMInstance5.PWMPulseWidthCountZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38547),
            .ce(N__19652),
            .sr(N__35737));
    defparam RST_ibuf_RNIUR47_LC_7_1_4.C_ON=1'b0;
    defparam RST_ibuf_RNIUR47_LC_7_1_4.SEQ_MODE=4'b0000;
    defparam RST_ibuf_RNIUR47_LC_7_1_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 RST_ibuf_RNIUR47_LC_7_1_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34515),
            .lcout(RST_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.delayedCh_B_0_LC_7_1_5 .C_ON=1'b0;
    defparam \QuadInstance0.delayedCh_B_0_LC_7_1_5 .SEQ_MODE=4'b1000;
    defparam \QuadInstance0.delayedCh_B_0_LC_7_1_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance0.delayedCh_B_0_LC_7_1_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15201),
            .lcout(\QuadInstance0.delayedCh_BZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38670),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance1.periodCounter_RNIFA3I1_3_LC_7_2_0 .C_ON=1'b0;
    defparam \PWMInstance1.periodCounter_RNIFA3I1_3_LC_7_2_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance1.periodCounter_RNIFA3I1_3_LC_7_2_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \PWMInstance1.periodCounter_RNIFA3I1_3_LC_7_2_0  (
            .in0(N__16201),
            .in1(N__16129),
            .in2(N__16349),
            .in3(N__16240),
            .lcout(\PWMInstance1.un1_periodCounter12_1_0_a2_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_7_2_1 .C_ON=1'b0;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_7_2_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_7_2_1 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \PWMInstance1.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_7_2_1  (
            .in0(N__16022),
            .in1(N__15312),
            .in2(N__16242),
            .in3(N__15318),
            .lcout(\PWMInstance1.un1_PWMPulseWidthCount_0_I_9_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance1.PWMPulseWidthCount_esr_2_LC_7_2_2 .C_ON=1'b0;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_2_LC_7_2_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_2_LC_7_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance1.PWMPulseWidthCount_esr_2_LC_7_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31608),
            .lcout(\PWMInstance1.PWMPulseWidthCountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38658),
            .ce(N__16827),
            .sr(N__35676));
    defparam \PWMInstance1.PWMPulseWidthCount_esr_3_LC_7_2_3 .C_ON=1'b0;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_3_LC_7_2_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_3_LC_7_2_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance1.PWMPulseWidthCount_esr_3_LC_7_2_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32091),
            .lcout(\PWMInstance1.PWMPulseWidthCountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38658),
            .ce(N__16827),
            .sr(N__35676));
    defparam \PWMInstance1.periodCounter_RNIT6VP_2_LC_7_2_4 .C_ON=1'b0;
    defparam \PWMInstance1.periodCounter_RNIT6VP_2_LC_7_2_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance1.periodCounter_RNIT6VP_2_LC_7_2_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \PWMInstance1.periodCounter_RNIT6VP_2_LC_7_2_4  (
            .in0(_gnd_net_),
            .in1(N__16267),
            .in2(_gnd_net_),
            .in3(N__16021),
            .lcout(),
            .ltout(\PWMInstance1.un1_periodCounter12_1_0_a2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance1.periodCounter_RNIUIR12_4_LC_7_2_5 .C_ON=1'b0;
    defparam \PWMInstance1.periodCounter_RNIUIR12_4_LC_7_2_5 .SEQ_MODE=4'b0000;
    defparam \PWMInstance1.periodCounter_RNIUIR12_4_LC_7_2_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \PWMInstance1.periodCounter_RNIUIR12_4_LC_7_2_5  (
            .in0(N__16318),
            .in1(N__16102),
            .in2(N__15303),
            .in3(N__16220),
            .lcout(\PWMInstance1.un1_periodCounter12_1_0_a2_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_7_2_6 .C_ON=1'b0;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_7_2_6 .SEQ_MODE=4'b0000;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_7_2_6 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \PWMInstance1.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_7_2_6  (
            .in0(N__16219),
            .in1(N__15354),
            .in2(N__16203),
            .in3(N__15300),
            .lcout(\PWMInstance1.un1_PWMPulseWidthCount_0_I_15_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance1.PWMPulseWidthCount_esr_4_LC_7_2_7 .C_ON=1'b0;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_4_LC_7_2_7 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_4_LC_7_2_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \PWMInstance1.PWMPulseWidthCount_esr_4_LC_7_2_7  (
            .in0(N__36525),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PWMInstance1.PWMPulseWidthCountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38658),
            .ce(N__16827),
            .sr(N__35676));
    defparam \PWMInstance1.periodCounter_RNIE93I1_0_LC_7_3_0 .C_ON=1'b0;
    defparam \PWMInstance1.periodCounter_RNIE93I1_0_LC_7_3_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance1.periodCounter_RNIE93I1_0_LC_7_3_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \PWMInstance1.periodCounter_RNIE93I1_0_LC_7_3_0  (
            .in0(N__16044),
            .in1(N__16295),
            .in2(N__16182),
            .in3(N__16151),
            .lcout(\PWMInstance1.un1_periodCounter12_1_0_a2_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_7_3_1 .C_ON=1'b0;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_7_3_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_7_3_1 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \PWMInstance1.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_7_3_1  (
            .in0(N__15387),
            .in1(N__16043),
            .in2(N__15396),
            .in3(N__16619),
            .lcout(\PWMInstance1.un1_PWMPulseWidthCount_0_I_1_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance1.PWMPulseWidthCount_esr_0_LC_7_3_2 .C_ON=1'b0;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_0_LC_7_3_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_0_LC_7_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance1.PWMPulseWidthCount_esr_0_LC_7_3_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31435),
            .lcout(\PWMInstance1.PWMPulseWidthCountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38648),
            .ce(N__16823),
            .sr(N__35677));
    defparam \PWMInstance1.PWMPulseWidthCount_esr_1_LC_7_3_3 .C_ON=1'b0;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_1_LC_7_3_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_1_LC_7_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance1.PWMPulseWidthCount_esr_1_LC_7_3_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31279),
            .lcout(\PWMInstance1.PWMPulseWidthCountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38648),
            .ce(N__16823),
            .sr(N__35677));
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_7_3_4 .C_ON=1'b0;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_7_3_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_7_3_4 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \PWMInstance1.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_7_3_4  (
            .in0(N__16178),
            .in1(N__15336),
            .in2(N__15381),
            .in3(N__16682),
            .lcout(\PWMInstance1.un1_PWMPulseWidthCount_0_I_27_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_7_3_7 .C_ON=1'b0;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_7_3_7 .SEQ_MODE=4'b0000;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_7_3_7 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance1.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_7_3_7  (
            .in0(N__15345),
            .in1(N__16150),
            .in2(N__16131),
            .in3(N__15366),
            .lcout(\PWMInstance1.un1_PWMPulseWidthCount_0_I_45_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance1.PWMPulseWidthCount_esr_13_LC_7_4_0 .C_ON=1'b0;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_13_LC_7_4_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_13_LC_7_4_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \PWMInstance1.PWMPulseWidthCount_esr_13_LC_7_4_0  (
            .in0(N__28728),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PWMInstance1.PWMPulseWidthCountZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38638),
            .ce(N__16825),
            .sr(N__35679));
    defparam \PWMInstance1.PWMPulseWidthCount_esr_5_LC_7_4_1 .C_ON=1'b0;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_5_LC_7_4_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_5_LC_7_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance1.PWMPulseWidthCount_esr_5_LC_7_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36377),
            .lcout(\PWMInstance1.PWMPulseWidthCountZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38638),
            .ce(N__16825),
            .sr(N__35679));
    defparam \PWMInstance1.PWMPulseWidthCount_esr_9_LC_7_4_3 .C_ON=1'b0;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_9_LC_7_4_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_9_LC_7_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance1.PWMPulseWidthCount_esr_9_LC_7_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28584),
            .lcout(\PWMInstance1.PWMPulseWidthCountZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38638),
            .ce(N__16825),
            .sr(N__35679));
    defparam \PWMInstance1.PWMPulseWidthCount_esr_6_LC_7_4_5 .C_ON=1'b0;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_6_LC_7_4_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_6_LC_7_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance1.PWMPulseWidthCount_esr_6_LC_7_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31124),
            .lcout(\PWMInstance1.PWMPulseWidthCountZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38638),
            .ce(N__16825),
            .sr(N__35679));
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_7_5_0 .C_ON=1'b0;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_7_5_0 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance1.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_7_5_0  (
            .in0(N__15438),
            .in1(N__15330),
            .in2(N__16659),
            .in3(N__16272),
            .lcout(\PWMInstance1.un1_PWMPulseWidthCount_0_I_21_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance1.PWMPulseWidthCount_esr_15_LC_7_5_2 .C_ON=1'b0;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_15_LC_7_5_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_15_LC_7_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance1.PWMPulseWidthCount_esr_15_LC_7_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31918),
            .lcout(\PWMInstance1.PWMPulseWidthCountZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38627),
            .ce(N__16824),
            .sr(N__35680));
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_7_5_3 .C_ON=1'b0;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_7_5_3 .SEQ_MODE=4'b0000;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_7_5_3 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \PWMInstance1.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_7_5_3  (
            .in0(N__16107),
            .in1(N__16365),
            .in2(N__15432),
            .in3(N__16350),
            .lcout(\PWMInstance1.un1_PWMPulseWidthCount_0_I_33_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_7_5_6 .C_ON=1'b0;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_7_5_6 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance1.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_7_5_6  (
            .in0(N__16323),
            .in1(N__16299),
            .in2(N__16374),
            .in3(N__15417),
            .lcout(\PWMInstance1.un1_PWMPulseWidthCount_0_I_39_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.un1_Quad_cry_0_c_LC_7_6_0 .C_ON=1'b1;
    defparam \QuadInstance2.un1_Quad_cry_0_c_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.un1_Quad_cry_0_c_LC_7_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \QuadInstance2.un1_Quad_cry_0_c_LC_7_6_0  (
            .in0(_gnd_net_),
            .in1(N__18529),
            .in2(N__30845),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_6_0_),
            .carryout(\QuadInstance2.un1_Quad_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_RNO_0_1_LC_7_6_1 .C_ON=1'b1;
    defparam \QuadInstance2.Quad_RNO_0_1_LC_7_6_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNO_0_1_LC_7_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance2.Quad_RNO_0_1_LC_7_6_1  (
            .in0(_gnd_net_),
            .in1(N__23834),
            .in2(N__15528),
            .in3(N__15411),
            .lcout(\QuadInstance2.Quad_RNO_0_1_1 ),
            .ltout(),
            .carryin(\QuadInstance2.un1_Quad_cry_0 ),
            .carryout(\QuadInstance2.un1_Quad_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_RNO_0_2_LC_7_6_2 .C_ON=1'b1;
    defparam \QuadInstance2.Quad_RNO_0_2_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNO_0_2_LC_7_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance2.Quad_RNO_0_2_LC_7_6_2  (
            .in0(_gnd_net_),
            .in1(N__30461),
            .in2(N__15627),
            .in3(N__15408),
            .lcout(\QuadInstance2.Quad_RNO_0_2_2 ),
            .ltout(),
            .carryin(\QuadInstance2.un1_Quad_cry_1 ),
            .carryout(\QuadInstance2.un1_Quad_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_RNO_0_3_LC_7_6_3 .C_ON=1'b1;
    defparam \QuadInstance2.Quad_RNO_0_3_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNO_0_3_LC_7_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance2.Quad_RNO_0_3_LC_7_6_3  (
            .in0(_gnd_net_),
            .in1(N__24406),
            .in2(N__15612),
            .in3(N__15405),
            .lcout(\QuadInstance2.Quad_RNO_0_2_3 ),
            .ltout(),
            .carryin(\QuadInstance2.un1_Quad_cry_2 ),
            .carryout(\QuadInstance2.un1_Quad_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_RNO_0_4_LC_7_6_4 .C_ON=1'b1;
    defparam \QuadInstance2.Quad_RNO_0_4_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNO_0_4_LC_7_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance2.Quad_RNO_0_4_LC_7_6_4  (
            .in0(_gnd_net_),
            .in1(N__21296),
            .in2(N__15477),
            .in3(N__15402),
            .lcout(\QuadInstance2.Quad_RNO_0_2_4 ),
            .ltout(),
            .carryin(\QuadInstance2.un1_Quad_cry_3 ),
            .carryout(\QuadInstance2.un1_Quad_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_RNO_0_5_LC_7_6_5 .C_ON=1'b1;
    defparam \QuadInstance2.Quad_RNO_0_5_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNO_0_5_LC_7_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance2.Quad_RNO_0_5_LC_7_6_5  (
            .in0(_gnd_net_),
            .in1(N__23717),
            .in2(N__15600),
            .in3(N__15399),
            .lcout(\QuadInstance2.Quad_RNO_0_2_5 ),
            .ltout(),
            .carryin(\QuadInstance2.un1_Quad_cry_4 ),
            .carryout(\QuadInstance2.un1_Quad_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_RNO_0_6_LC_7_6_6 .C_ON=1'b1;
    defparam \QuadInstance2.Quad_RNO_0_6_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNO_0_6_LC_7_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance2.Quad_RNO_0_6_LC_7_6_6  (
            .in0(_gnd_net_),
            .in1(N__28300),
            .in2(N__15588),
            .in3(N__15465),
            .lcout(\QuadInstance2.Quad_RNO_0_2_6 ),
            .ltout(),
            .carryin(\QuadInstance2.un1_Quad_cry_5 ),
            .carryout(\QuadInstance2.un1_Quad_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_RNO_0_7_LC_7_6_7 .C_ON=1'b1;
    defparam \QuadInstance2.Quad_RNO_0_7_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNO_0_7_LC_7_6_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance2.Quad_RNO_0_7_LC_7_6_7  (
            .in0(_gnd_net_),
            .in1(N__26374),
            .in2(N__15498),
            .in3(N__15462),
            .lcout(\QuadInstance2.Quad_RNO_0_2_7 ),
            .ltout(),
            .carryin(\QuadInstance2.un1_Quad_cry_6 ),
            .carryout(\QuadInstance2.un1_Quad_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_RNO_0_8_LC_7_7_0 .C_ON=1'b1;
    defparam \QuadInstance2.Quad_RNO_0_8_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNO_0_8_LC_7_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance2.Quad_RNO_0_8_LC_7_7_0  (
            .in0(_gnd_net_),
            .in1(N__30703),
            .in2(N__15486),
            .in3(N__15459),
            .lcout(\QuadInstance2.Quad_RNO_0_2_8 ),
            .ltout(),
            .carryin(bfn_7_7_0_),
            .carryout(\QuadInstance2.un1_Quad_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_RNO_0_9_LC_7_7_1 .C_ON=1'b1;
    defparam \QuadInstance2.Quad_RNO_0_9_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNO_0_9_LC_7_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance2.Quad_RNO_0_9_LC_7_7_1  (
            .in0(_gnd_net_),
            .in1(N__25438),
            .in2(N__15546),
            .in3(N__15456),
            .lcout(\QuadInstance2.Quad_RNO_0_2_9 ),
            .ltout(),
            .carryin(\QuadInstance2.un1_Quad_cry_8 ),
            .carryout(\QuadInstance2.un1_Quad_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_RNO_0_10_LC_7_7_2 .C_ON=1'b1;
    defparam \QuadInstance2.Quad_RNO_0_10_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNO_0_10_LC_7_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance2.Quad_RNO_0_10_LC_7_7_2  (
            .in0(_gnd_net_),
            .in1(N__34675),
            .in2(N__15516),
            .in3(N__15453),
            .lcout(\QuadInstance2.Quad_RNO_0_2_10 ),
            .ltout(),
            .carryin(\QuadInstance2.un1_Quad_cry_9 ),
            .carryout(\QuadInstance2.un1_Quad_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_RNO_0_11_LC_7_7_3 .C_ON=1'b1;
    defparam \QuadInstance2.Quad_RNO_0_11_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNO_0_11_LC_7_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance2.Quad_RNO_0_11_LC_7_7_3  (
            .in0(_gnd_net_),
            .in1(N__22451),
            .in2(N__15537),
            .in3(N__15450),
            .lcout(\QuadInstance2.Quad_RNO_0_2_11 ),
            .ltout(),
            .carryin(\QuadInstance2.un1_Quad_cry_10 ),
            .carryout(\QuadInstance2.un1_Quad_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_RNO_0_12_LC_7_7_4 .C_ON=1'b1;
    defparam \QuadInstance2.Quad_RNO_0_12_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNO_0_12_LC_7_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance2.Quad_RNO_0_12_LC_7_7_4  (
            .in0(_gnd_net_),
            .in1(N__22351),
            .in2(N__15507),
            .in3(N__15447),
            .lcout(\QuadInstance2.Quad_RNO_0_2_12 ),
            .ltout(),
            .carryin(\QuadInstance2.un1_Quad_cry_11 ),
            .carryout(\QuadInstance2.un1_Quad_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_RNO_0_13_LC_7_7_5 .C_ON=1'b1;
    defparam \QuadInstance2.Quad_RNO_0_13_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNO_0_13_LC_7_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance2.Quad_RNO_0_13_LC_7_7_5  (
            .in0(_gnd_net_),
            .in1(N__19973),
            .in2(N__17520),
            .in3(N__15444),
            .lcout(\QuadInstance2.Quad_RNO_0_2_13 ),
            .ltout(),
            .carryin(\QuadInstance2.un1_Quad_cry_12 ),
            .carryout(\QuadInstance2.un1_Quad_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_RNO_0_14_LC_7_7_6 .C_ON=1'b1;
    defparam \QuadInstance2.Quad_RNO_0_14_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNO_0_14_LC_7_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance2.Quad_RNO_0_14_LC_7_7_6  (
            .in0(_gnd_net_),
            .in1(N__15714),
            .in2(N__20047),
            .in3(N__15441),
            .lcout(\QuadInstance2.Quad_RNO_0_2_14 ),
            .ltout(),
            .carryin(\QuadInstance2.un1_Quad_cry_13 ),
            .carryout(\QuadInstance2.un1_Quad_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_15_LC_7_7_7 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_15_LC_7_7_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance2.Quad_15_LC_7_7_7 .LUT_INIT=16'b1101000111100010;
    LogicCell40 \QuadInstance2.Quad_15_LC_7_7_7  (
            .in0(N__15639),
            .in1(N__22159),
            .in2(N__31923),
            .in3(N__15549),
            .lcout(dataRead2_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38606),
            .ce(),
            .sr(N__35684));
    defparam \QuadInstance2.Quad_RNI8TLE2_9_LC_7_8_0 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_RNI8TLE2_9_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNI8TLE2_9_LC_7_8_0 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance2.Quad_RNI8TLE2_9_LC_7_8_0  (
            .in0(N__25442),
            .in1(N__22102),
            .in2(N__18518),
            .in3(N__17572),
            .lcout(\QuadInstance2.Quad_RNI8TLE2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_RNIHU2G2_11_LC_7_8_1 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_RNIHU2G2_11_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNIHU2G2_11_LC_7_8_1 .LUT_INIT=16'b1010111100000000;
    LogicCell40 \QuadInstance2.Quad_RNIHU2G2_11_LC_7_8_1  (
            .in0(N__22105),
            .in1(N__22455),
            .in2(N__17592),
            .in3(N__18503),
            .lcout(\QuadInstance2.Quad_RNIHU2G2Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_RNI0LLE2_1_LC_7_8_2 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_RNI0LLE2_1_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNI0LLE2_1_LC_7_8_2 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance2.Quad_RNI0LLE2_1_LC_7_8_2  (
            .in0(N__23835),
            .in1(N__22098),
            .in2(N__18516),
            .in3(N__17561),
            .lcout(\QuadInstance2.Quad_RNI0LLE2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_RNIGT2G2_10_LC_7_8_3 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_RNIGT2G2_10_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNIGT2G2_10_LC_7_8_3 .LUT_INIT=16'b1010111100000000;
    LogicCell40 \QuadInstance2.Quad_RNIGT2G2_10_LC_7_8_3  (
            .in0(N__22103),
            .in1(N__34676),
            .in2(N__17591),
            .in3(N__18499),
            .lcout(\QuadInstance2.Quad_RNIGT2G2Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_RNIIV2G2_12_LC_7_8_4 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_RNIIV2G2_12_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNIIV2G2_12_LC_7_8_4 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance2.Quad_RNIIV2G2_12_LC_7_8_4  (
            .in0(N__22352),
            .in1(N__22104),
            .in2(N__18519),
            .in3(N__17576),
            .lcout(\QuadInstance2.Quad_RNIIV2G2Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_RNI6RLE2_7_LC_7_8_5 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_RNI6RLE2_7_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNI6RLE2_7_LC_7_8_5 .LUT_INIT=16'b1010111100000000;
    LogicCell40 \QuadInstance2.Quad_RNI6RLE2_7_LC_7_8_5  (
            .in0(N__22100),
            .in1(N__26375),
            .in2(N__17590),
            .in3(N__18492),
            .lcout(\QuadInstance2.Quad_RNI6RLE2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_RNI7SLE2_8_LC_7_8_6 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_RNI7SLE2_8_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNI7SLE2_8_LC_7_8_6 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance2.Quad_RNI7SLE2_8_LC_7_8_6  (
            .in0(N__30711),
            .in1(N__22101),
            .in2(N__18517),
            .in3(N__17568),
            .lcout(\QuadInstance2.Quad_RNI7SLE2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_RNI3OLE2_4_LC_7_8_7 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_RNI3OLE2_4_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNI3OLE2_4_LC_7_8_7 .LUT_INIT=16'b1010111100000000;
    LogicCell40 \QuadInstance2.Quad_RNI3OLE2_4_LC_7_8_7  (
            .in0(N__22099),
            .in1(N__21297),
            .in2(N__17589),
            .in3(N__18491),
            .lcout(\QuadInstance2.Quad_RNI3OLE2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_RNO_0_15_LC_7_9_0 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_RNO_0_15_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNO_0_15_LC_7_9_0 .LUT_INIT=16'b0100101111110000;
    LogicCell40 \QuadInstance2.Quad_RNO_0_15_LC_7_9_0  (
            .in0(N__22110),
            .in1(N__17584),
            .in2(N__24314),
            .in3(N__18507),
            .lcout(\QuadInstance2.un1_Quad_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.delayedCh_A_RNIK9UB1_2_LC_7_9_1 .C_ON=1'b0;
    defparam \QuadInstance2.delayedCh_A_RNIK9UB1_2_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.delayedCh_A_RNIK9UB1_2_LC_7_9_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \QuadInstance2.delayedCh_A_RNIK9UB1_2_LC_7_9_1  (
            .in0(N__15555),
            .in1(N__15693),
            .in2(N__15575),
            .in3(N__15704),
            .lcout(\QuadInstance2.count_enable ),
            .ltout(\QuadInstance2.count_enable_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_RNI1MLE2_2_LC_7_9_2 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_RNI1MLE2_2_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNI1MLE2_2_LC_7_9_2 .LUT_INIT=16'b1010000011110000;
    LogicCell40 \QuadInstance2.Quad_RNI1MLE2_2_LC_7_9_2  (
            .in0(N__22106),
            .in1(N__30465),
            .in2(N__15630),
            .in3(N__17577),
            .lcout(\QuadInstance2.Quad_RNI1MLE2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.delayedCh_B_RNIO04T_2_LC_7_9_3 .C_ON=1'b0;
    defparam \QuadInstance2.delayedCh_B_RNIO04T_2_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.delayedCh_B_RNIO04T_2_LC_7_9_3 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \QuadInstance2.delayedCh_B_RNIO04T_2_LC_7_9_3  (
            .in0(N__34471),
            .in1(_gnd_net_),
            .in2(N__15576),
            .in3(N__15692),
            .lcout(\QuadInstance2.un1_count_enable_i_a2_0_1 ),
            .ltout(\QuadInstance2.un1_count_enable_i_a2_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_RNI2NLE2_3_LC_7_9_4 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_RNI2NLE2_3_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNI2NLE2_3_LC_7_9_4 .LUT_INIT=16'b1010111100000000;
    LogicCell40 \QuadInstance2.Quad_RNI2NLE2_3_LC_7_9_4  (
            .in0(N__22107),
            .in1(N__24414),
            .in2(N__15615),
            .in3(N__18504),
            .lcout(\QuadInstance2.Quad_RNI2NLE2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_RNI4PLE2_5_LC_7_9_5 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_RNI4PLE2_5_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNI4PLE2_5_LC_7_9_5 .LUT_INIT=16'b1000101010001010;
    LogicCell40 \QuadInstance2.Quad_RNI4PLE2_5_LC_7_9_5  (
            .in0(N__18506),
            .in1(N__22109),
            .in2(N__17594),
            .in3(N__23718),
            .lcout(\QuadInstance2.Quad_RNI4PLE2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNO_0_15_LC_7_9_6 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_RNO_0_15_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNO_0_15_LC_7_9_6 .LUT_INIT=16'b0011100111001100;
    LogicCell40 \QuadInstance7.Quad_RNO_0_15_LC_7_9_6  (
            .in0(N__16522),
            .in1(N__24290),
            .in2(N__26011),
            .in3(N__21795),
            .lcout(\QuadInstance7.un1_Quad_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_RNI5QLE2_6_LC_7_9_7 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_RNI5QLE2_6_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNI5QLE2_6_LC_7_9_7 .LUT_INIT=16'b1000101010001010;
    LogicCell40 \QuadInstance2.Quad_RNI5QLE2_6_LC_7_9_7  (
            .in0(N__18505),
            .in1(N__22108),
            .in2(N__17593),
            .in3(N__28305),
            .lcout(\QuadInstance2.Quad_RNI5QLE2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.delayedCh_A_1_LC_7_10_0 .C_ON=1'b0;
    defparam \QuadInstance2.delayedCh_A_1_LC_7_10_0 .SEQ_MODE=4'b1000;
    defparam \QuadInstance2.delayedCh_A_1_LC_7_10_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \QuadInstance2.delayedCh_A_1_LC_7_10_0  (
            .in0(N__21339),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\QuadInstance2.delayedCh_AZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38575),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.delayedCh_A_2_LC_7_10_2 .C_ON=1'b0;
    defparam \QuadInstance2.delayedCh_A_2_LC_7_10_2 .SEQ_MODE=4'b1000;
    defparam \QuadInstance2.delayedCh_A_2_LC_7_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance2.delayedCh_A_2_LC_7_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15574),
            .lcout(\QuadInstance2.delayedCh_AZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38575),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.delayedCh_B_1_LC_7_10_3 .C_ON=1'b0;
    defparam \QuadInstance2.delayedCh_B_1_LC_7_10_3 .SEQ_MODE=4'b1000;
    defparam \QuadInstance2.delayedCh_B_1_LC_7_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance2.delayedCh_B_1_LC_7_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23313),
            .lcout(\QuadInstance2.delayedCh_BZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38575),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_RNIK13G2_14_LC_7_10_4 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_RNIK13G2_14_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNIK13G2_14_LC_7_10_4 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \QuadInstance2.Quad_RNIK13G2_14_LC_7_10_4  (
            .in0(N__22150),
            .in1(N__18515),
            .in2(N__20049),
            .in3(N__17588),
            .lcout(\QuadInstance2.Quad_RNIK13G2Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.delayedCh_B_2_LC_7_10_5 .C_ON=1'b0;
    defparam \QuadInstance2.delayedCh_B_2_LC_7_10_5 .SEQ_MODE=4'b1000;
    defparam \QuadInstance2.delayedCh_B_2_LC_7_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance2.delayedCh_B_2_LC_7_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15705),
            .lcout(\QuadInstance2.delayedCh_BZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38575),
            .ce(),
            .sr(_gnd_net_));
    defparam pwmWrite_fast_0_LC_7_10_6.C_ON=1'b0;
    defparam pwmWrite_fast_0_LC_7_10_6.SEQ_MODE=4'b1000;
    defparam pwmWrite_fast_0_LC_7_10_6.LUT_INIT=16'b0000000100000000;
    LogicCell40 pwmWrite_fast_0_LC_7_10_6 (
            .in0(N__33846),
            .in1(N__33659),
            .in2(N__33441),
            .in3(N__33231),
            .lcout(pwmWrite_fastZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38575),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_1_c_LC_7_11_0 .C_ON=1'b1;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_1_c_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_1_c_LC_7_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance1.un1_PWMPulseWidthCount_0_I_1_c_LC_7_11_0  (
            .in0(_gnd_net_),
            .in1(N__15684),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_11_0_),
            .carryout(\PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_9_c_LC_7_11_1 .C_ON=1'b1;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_9_c_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_9_c_LC_7_11_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance1.un1_PWMPulseWidthCount_0_I_9_c_LC_7_11_1  (
            .in0(_gnd_net_),
            .in1(N__15675),
            .in2(N__32472),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_0 ),
            .carryout(\PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_15_c_LC_7_11_2 .C_ON=1'b1;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_15_c_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_15_c_LC_7_11_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance1.un1_PWMPulseWidthCount_0_I_15_c_LC_7_11_2  (
            .in0(_gnd_net_),
            .in1(N__15666),
            .in2(N__32466),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_1 ),
            .carryout(\PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_27_c_LC_7_11_3 .C_ON=1'b1;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_27_c_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_27_c_LC_7_11_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance1.un1_PWMPulseWidthCount_0_I_27_c_LC_7_11_3  (
            .in0(_gnd_net_),
            .in1(N__15651),
            .in2(N__32470),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_2 ),
            .carryout(\PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_45_c_LC_7_11_4 .C_ON=1'b1;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_45_c_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_45_c_LC_7_11_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance1.un1_PWMPulseWidthCount_0_I_45_c_LC_7_11_4  (
            .in0(_gnd_net_),
            .in1(N__15783),
            .in2(N__32468),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_3 ),
            .carryout(\PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_33_c_LC_7_11_5 .C_ON=1'b1;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_33_c_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_33_c_LC_7_11_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance1.un1_PWMPulseWidthCount_0_I_33_c_LC_7_11_5  (
            .in0(_gnd_net_),
            .in1(N__15771),
            .in2(N__32471),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_4 ),
            .carryout(\PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_39_c_LC_7_11_6 .C_ON=1'b1;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_39_c_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_39_c_LC_7_11_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance1.un1_PWMPulseWidthCount_0_I_39_c_LC_7_11_6  (
            .in0(_gnd_net_),
            .in1(N__15759),
            .in2(N__32467),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_5 ),
            .carryout(\PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_21_c_LC_7_11_7 .C_ON=1'b1;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_21_c_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \PWMInstance1.un1_PWMPulseWidthCount_0_I_21_c_LC_7_11_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance1.un1_PWMPulseWidthCount_0_I_21_c_LC_7_11_7  (
            .in0(_gnd_net_),
            .in1(N__15747),
            .in2(N__32469),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_6 ),
            .carryout(\PWMInstance1.un1_PWMPulseWidthCount_0_data_tmp_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance1.out_LC_7_12_0 .C_ON=1'b0;
    defparam \PWMInstance1.out_LC_7_12_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.out_LC_7_12_0 .LUT_INIT=16'b1111101011110010;
    LogicCell40 \PWMInstance1.out_LC_7_12_0  (
            .in0(N__15725),
            .in1(N__16833),
            .in2(N__16999),
            .in3(N__15738),
            .lcout(PWM1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38559),
            .ce(),
            .sr(N__35719));
    defparam \PWMInstance0.PWMPulseWidthCount_esr_13_LC_7_13_0 .C_ON=1'b0;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_13_LC_7_13_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_13_LC_7_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance0.PWMPulseWidthCount_esr_13_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28723),
            .lcout(\PWMInstance0.PWMPulseWidthCountZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38552),
            .ce(N__18233),
            .sr(N__35727));
    defparam \PWMInstance0.PWMPulseWidthCount_esr_5_LC_7_13_1 .C_ON=1'b0;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_5_LC_7_13_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_5_LC_7_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance0.PWMPulseWidthCount_esr_5_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36367),
            .lcout(\PWMInstance0.PWMPulseWidthCountZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38552),
            .ce(N__18233),
            .sr(N__35727));
    defparam \PWMInstance0.PWMPulseWidthCount_esr_8_LC_7_13_2 .C_ON=1'b0;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_8_LC_7_13_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_8_LC_7_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance0.PWMPulseWidthCount_esr_8_LC_7_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28992),
            .lcout(\PWMInstance0.PWMPulseWidthCountZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38552),
            .ce(N__18233),
            .sr(N__35727));
    defparam \PWMInstance0.PWMPulseWidthCount_esr_9_LC_7_13_3 .C_ON=1'b0;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_9_LC_7_13_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_9_LC_7_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance0.PWMPulseWidthCount_esr_9_LC_7_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28576),
            .lcout(\PWMInstance0.PWMPulseWidthCountZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38552),
            .ce(N__18233),
            .sr(N__35727));
    defparam \PWMInstance0.PWMPulseWidthCount_esr_12_LC_7_13_5 .C_ON=1'b0;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_12_LC_7_13_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_12_LC_7_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance0.PWMPulseWidthCount_esr_12_LC_7_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28870),
            .lcout(\PWMInstance0.PWMPulseWidthCountZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38552),
            .ce(N__18233),
            .sr(N__35727));
    defparam \PWMInstance0.PWMPulseWidthCount_esr_6_LC_7_13_6 .C_ON=1'b0;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_6_LC_7_13_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_6_LC_7_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance0.PWMPulseWidthCount_esr_6_LC_7_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31114),
            .lcout(\PWMInstance0.PWMPulseWidthCountZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38552),
            .ce(N__18233),
            .sr(N__35727));
    defparam \PWMInstance0.PWMPulseWidthCount_esr_4_LC_7_13_7 .C_ON=1'b0;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_4_LC_7_13_7 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_4_LC_7_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance0.PWMPulseWidthCount_esr_4_LC_7_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36513),
            .lcout(\PWMInstance0.PWMPulseWidthCountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38552),
            .ce(N__18233),
            .sr(N__35727));
    defparam \PWMInstance0.periodCounter_RNIB5GO1_11_LC_7_14_0 .C_ON=1'b0;
    defparam \PWMInstance0.periodCounter_RNIB5GO1_11_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance0.periodCounter_RNIB5GO1_11_LC_7_14_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \PWMInstance0.periodCounter_RNIB5GO1_11_LC_7_14_0  (
            .in0(N__15938),
            .in1(N__16904),
            .in2(N__17088),
            .in3(N__15983),
            .lcout(\PWMInstance0.un1_periodCounter12_1_0_a2_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_7_14_1 .C_ON=1'b0;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_7_14_1 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \PWMInstance0.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_7_14_1  (
            .in0(N__16005),
            .in1(N__15807),
            .in2(N__15984),
            .in3(N__15813),
            .lcout(\PWMInstance0.un1_PWMPulseWidthCount_0_I_9_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance0.PWMPulseWidthCount_esr_2_LC_7_14_2 .C_ON=1'b0;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_2_LC_7_14_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_2_LC_7_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance0.PWMPulseWidthCount_esr_2_LC_7_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31603),
            .lcout(\PWMInstance0.PWMPulseWidthCountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38548),
            .ce(N__18235),
            .sr(N__35738));
    defparam \PWMInstance0.PWMPulseWidthCount_esr_3_LC_7_14_3 .C_ON=1'b0;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_3_LC_7_14_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_3_LC_7_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance0.PWMPulseWidthCount_esr_3_LC_7_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32082),
            .lcout(\PWMInstance0.PWMPulseWidthCountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38548),
            .ce(N__18235),
            .sr(N__35738));
    defparam \PWMInstance0.periodCounter_RNIR3TO_14_LC_7_14_4 .C_ON=1'b0;
    defparam \PWMInstance0.periodCounter_RNIR3TO_14_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance0.periodCounter_RNIR3TO_14_LC_7_14_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \PWMInstance0.periodCounter_RNIR3TO_14_LC_7_14_4  (
            .in0(_gnd_net_),
            .in1(N__17147),
            .in2(_gnd_net_),
            .in3(N__16004),
            .lcout(),
            .ltout(\PWMInstance0.un1_periodCounter12_1_0_a2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance0.periodCounter_RNIPQTQ1_10_LC_7_14_5 .C_ON=1'b0;
    defparam \PWMInstance0.periodCounter_RNIPQTQ1_10_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \PWMInstance0.periodCounter_RNIPQTQ1_10_LC_7_14_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \PWMInstance0.periodCounter_RNIPQTQ1_10_LC_7_14_5  (
            .in0(N__15960),
            .in1(N__17027),
            .in2(N__15798),
            .in3(N__17112),
            .lcout(\PWMInstance0.un1_periodCounter12_1_0_a2_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_7_14_6 .C_ON=1'b0;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_7_14_6 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance0.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_7_14_6  (
            .in0(N__15795),
            .in1(N__15959),
            .in2(N__15939),
            .in3(N__15789),
            .lcout(\PWMInstance0.un1_PWMPulseWidthCount_0_I_15_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance0.out_RNO_0_LC_7_15_0 .C_ON=1'b0;
    defparam \PWMInstance0.out_RNO_0_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance0.out_RNO_0_LC_7_15_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \PWMInstance0.out_RNO_0_LC_7_15_0  (
            .in0(N__15868),
            .in1(N__15900),
            .in2(N__15888),
            .in3(N__16062),
            .lcout(\PWMInstance0.un1_periodCounter12_1_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance0.clkCount_0_LC_7_15_1 .C_ON=1'b0;
    defparam \PWMInstance0.clkCount_0_LC_7_15_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.clkCount_0_LC_7_15_1 .LUT_INIT=16'b1010101000010001;
    LogicCell40 \PWMInstance0.clkCount_0_LC_7_15_1  (
            .in0(N__16874),
            .in1(N__15886),
            .in2(_gnd_net_),
            .in3(N__15869),
            .lcout(\PWMInstance0.clkCountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38545),
            .ce(),
            .sr(N__35742));
    defparam \PWMInstance0.clkCount_1_LC_7_15_3 .C_ON=1'b0;
    defparam \PWMInstance0.clkCount_1_LC_7_15_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.clkCount_1_LC_7_15_3 .LUT_INIT=16'b1001100110001000;
    LogicCell40 \PWMInstance0.clkCount_1_LC_7_15_3  (
            .in0(N__16875),
            .in1(N__15887),
            .in2(_gnd_net_),
            .in3(N__15870),
            .lcout(\PWMInstance0.clkCountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38545),
            .ce(),
            .sr(N__35742));
    defparam \PWMInstance0.periodCounter_RNI2BTO_16_LC_7_15_4 .C_ON=1'b0;
    defparam \PWMInstance0.periodCounter_RNI2BTO_16_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance0.periodCounter_RNI2BTO_16_LC_7_15_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \PWMInstance0.periodCounter_RNI2BTO_16_LC_7_15_4  (
            .in0(_gnd_net_),
            .in1(N__16061),
            .in2(_gnd_net_),
            .in3(N__17194),
            .lcout(\PWMInstance0.un1_periodCounter12_1_0_a2_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance0.clkCount_RNIPL0S_0_LC_7_15_5 .C_ON=1'b0;
    defparam \PWMInstance0.clkCount_RNIPL0S_0_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \PWMInstance0.clkCount_RNIPL0S_0_LC_7_15_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \PWMInstance0.clkCount_RNIPL0S_0_LC_7_15_5  (
            .in0(N__15899),
            .in1(N__15882),
            .in2(_gnd_net_),
            .in3(N__15867),
            .lcout(\PWMInstance0.periodCounter12 ),
            .ltout(\PWMInstance0.periodCounter12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance0.periodCounter_RNIM4RD2_15_LC_7_15_6 .C_ON=1'b0;
    defparam \PWMInstance0.periodCounter_RNIM4RD2_15_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \PWMInstance0.periodCounter_RNIM4RD2_15_LC_7_15_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \PWMInstance0.periodCounter_RNIM4RD2_15_LC_7_15_6  (
            .in0(N__17171),
            .in1(N__18007),
            .in2(N__15855),
            .in3(N__15852),
            .lcout(),
            .ltout(\PWMInstance0.un1_periodCounter12_1_0_a2_0_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance0.periodCounter_RNI49PP7_10_LC_7_15_7 .C_ON=1'b0;
    defparam \PWMInstance0.periodCounter_RNI49PP7_10_LC_7_15_7 .SEQ_MODE=4'b0000;
    defparam \PWMInstance0.periodCounter_RNI49PP7_10_LC_7_15_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \PWMInstance0.periodCounter_RNI49PP7_10_LC_7_15_7  (
            .in0(N__15846),
            .in1(N__18045),
            .in2(N__15840),
            .in3(N__15837),
            .lcout(\PWMInstance0.out_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance0.periodCounter_0_LC_7_16_0 .C_ON=1'b1;
    defparam \PWMInstance0.periodCounter_0_LC_7_16_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.periodCounter_0_LC_7_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance0.periodCounter_0_LC_7_16_0  (
            .in0(_gnd_net_),
            .in1(N__18034),
            .in2(N__15831),
            .in3(N__15830),
            .lcout(\PWMInstance0.periodCounterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_7_16_0_),
            .carryout(\PWMInstance0.un1_periodCounter_2_cry_0 ),
            .clk(N__38544),
            .ce(),
            .sr(N__35303));
    defparam \PWMInstance0.periodCounter_1_LC_7_16_1 .C_ON=1'b1;
    defparam \PWMInstance0.periodCounter_1_LC_7_16_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.periodCounter_1_LC_7_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance0.periodCounter_1_LC_7_16_1  (
            .in0(_gnd_net_),
            .in1(N__18011),
            .in2(_gnd_net_),
            .in3(N__15816),
            .lcout(\PWMInstance0.periodCounterZ0Z_1 ),
            .ltout(),
            .carryin(\PWMInstance0.un1_periodCounter_2_cry_0 ),
            .carryout(\PWMInstance0.un1_periodCounter_2_cry_1 ),
            .clk(N__38544),
            .ce(),
            .sr(N__35303));
    defparam \PWMInstance0.periodCounter_2_LC_7_16_2 .C_ON=1'b1;
    defparam \PWMInstance0.periodCounter_2_LC_7_16_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.periodCounter_2_LC_7_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance0.periodCounter_2_LC_7_16_2  (
            .in0(_gnd_net_),
            .in1(N__16003),
            .in2(_gnd_net_),
            .in3(N__15987),
            .lcout(\PWMInstance0.periodCounterZ0Z_2 ),
            .ltout(),
            .carryin(\PWMInstance0.un1_periodCounter_2_cry_1 ),
            .carryout(\PWMInstance0.un1_periodCounter_2_cry_2 ),
            .clk(N__38544),
            .ce(),
            .sr(N__35303));
    defparam \PWMInstance0.periodCounter_3_LC_7_16_3 .C_ON=1'b1;
    defparam \PWMInstance0.periodCounter_3_LC_7_16_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.periodCounter_3_LC_7_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance0.periodCounter_3_LC_7_16_3  (
            .in0(_gnd_net_),
            .in1(N__15979),
            .in2(_gnd_net_),
            .in3(N__15963),
            .lcout(\PWMInstance0.periodCounterZ0Z_3 ),
            .ltout(),
            .carryin(\PWMInstance0.un1_periodCounter_2_cry_2 ),
            .carryout(\PWMInstance0.un1_periodCounter_2_cry_3 ),
            .clk(N__38544),
            .ce(),
            .sr(N__35303));
    defparam \PWMInstance0.periodCounter_4_LC_7_16_4 .C_ON=1'b1;
    defparam \PWMInstance0.periodCounter_4_LC_7_16_4 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.periodCounter_4_LC_7_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance0.periodCounter_4_LC_7_16_4  (
            .in0(_gnd_net_),
            .in1(N__15958),
            .in2(_gnd_net_),
            .in3(N__15942),
            .lcout(\PWMInstance0.periodCounterZ0Z_4 ),
            .ltout(),
            .carryin(\PWMInstance0.un1_periodCounter_2_cry_3 ),
            .carryout(\PWMInstance0.un1_periodCounter_2_cry_4 ),
            .clk(N__38544),
            .ce(),
            .sr(N__35303));
    defparam \PWMInstance0.periodCounter_5_LC_7_16_5 .C_ON=1'b1;
    defparam \PWMInstance0.periodCounter_5_LC_7_16_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.periodCounter_5_LC_7_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance0.periodCounter_5_LC_7_16_5  (
            .in0(_gnd_net_),
            .in1(N__15934),
            .in2(_gnd_net_),
            .in3(N__15918),
            .lcout(\PWMInstance0.periodCounterZ0Z_5 ),
            .ltout(),
            .carryin(\PWMInstance0.un1_periodCounter_2_cry_4 ),
            .carryout(\PWMInstance0.un1_periodCounter_2_cry_5 ),
            .clk(N__38544),
            .ce(),
            .sr(N__35303));
    defparam \PWMInstance0.periodCounter_6_LC_7_16_6 .C_ON=1'b1;
    defparam \PWMInstance0.periodCounter_6_LC_7_16_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.periodCounter_6_LC_7_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance0.periodCounter_6_LC_7_16_6  (
            .in0(_gnd_net_),
            .in1(N__18100),
            .in2(_gnd_net_),
            .in3(N__15915),
            .lcout(\PWMInstance0.periodCounterZ0Z_6 ),
            .ltout(),
            .carryin(\PWMInstance0.un1_periodCounter_2_cry_5 ),
            .carryout(\PWMInstance0.un1_periodCounter_2_cry_6 ),
            .clk(N__38544),
            .ce(),
            .sr(N__35303));
    defparam \PWMInstance0.periodCounter_7_LC_7_16_7 .C_ON=1'b1;
    defparam \PWMInstance0.periodCounter_7_LC_7_16_7 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.periodCounter_7_LC_7_16_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance0.periodCounter_7_LC_7_16_7  (
            .in0(N__17284),
            .in1(N__17198),
            .in2(_gnd_net_),
            .in3(N__15912),
            .lcout(\PWMInstance0.periodCounterZ0Z_7 ),
            .ltout(),
            .carryin(\PWMInstance0.un1_periodCounter_2_cry_6 ),
            .carryout(\PWMInstance0.un1_periodCounter_2_cry_7 ),
            .clk(N__38544),
            .ce(),
            .sr(N__35303));
    defparam \PWMInstance0.periodCounter_8_LC_7_17_0 .C_ON=1'b1;
    defparam \PWMInstance0.periodCounter_8_LC_7_17_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.periodCounter_8_LC_7_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance0.periodCounter_8_LC_7_17_0  (
            .in0(_gnd_net_),
            .in1(N__18133),
            .in2(_gnd_net_),
            .in3(N__15909),
            .lcout(\PWMInstance0.periodCounterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_7_17_0_),
            .carryout(\PWMInstance0.un1_periodCounter_2_cry_8 ),
            .clk(N__38543),
            .ce(),
            .sr(N__35301));
    defparam \PWMInstance0.periodCounter_9_LC_7_17_1 .C_ON=1'b1;
    defparam \PWMInstance0.periodCounter_9_LC_7_17_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.periodCounter_9_LC_7_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance0.periodCounter_9_LC_7_17_1  (
            .in0(_gnd_net_),
            .in1(N__16900),
            .in2(_gnd_net_),
            .in3(N__15906),
            .lcout(\PWMInstance0.periodCounterZ0Z_9 ),
            .ltout(),
            .carryin(\PWMInstance0.un1_periodCounter_2_cry_8 ),
            .carryout(\PWMInstance0.un1_periodCounter_2_cry_9 ),
            .clk(N__38543),
            .ce(),
            .sr(N__35301));
    defparam \PWMInstance0.periodCounter_10_LC_7_17_2 .C_ON=1'b1;
    defparam \PWMInstance0.periodCounter_10_LC_7_17_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.periodCounter_10_LC_7_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance0.periodCounter_10_LC_7_17_2  (
            .in0(_gnd_net_),
            .in1(N__17110),
            .in2(_gnd_net_),
            .in3(N__15903),
            .lcout(\PWMInstance0.periodCounterZ0Z_10 ),
            .ltout(),
            .carryin(\PWMInstance0.un1_periodCounter_2_cry_9 ),
            .carryout(\PWMInstance0.un1_periodCounter_2_cry_10 ),
            .clk(N__38543),
            .ce(),
            .sr(N__35301));
    defparam \PWMInstance0.periodCounter_11_LC_7_17_3 .C_ON=1'b1;
    defparam \PWMInstance0.periodCounter_11_LC_7_17_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.periodCounter_11_LC_7_17_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance0.periodCounter_11_LC_7_17_3  (
            .in0(N__17289),
            .in1(N__17080),
            .in2(_gnd_net_),
            .in3(N__16080),
            .lcout(\PWMInstance0.periodCounterZ0Z_11 ),
            .ltout(),
            .carryin(\PWMInstance0.un1_periodCounter_2_cry_10 ),
            .carryout(\PWMInstance0.un1_periodCounter_2_cry_11 ),
            .clk(N__38543),
            .ce(),
            .sr(N__35301));
    defparam \PWMInstance0.periodCounter_12_LC_7_17_4 .C_ON=1'b1;
    defparam \PWMInstance0.periodCounter_12_LC_7_17_4 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.periodCounter_12_LC_7_17_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance0.periodCounter_12_LC_7_17_4  (
            .in0(N__17291),
            .in1(N__17026),
            .in2(_gnd_net_),
            .in3(N__16077),
            .lcout(\PWMInstance0.periodCounterZ0Z_12 ),
            .ltout(),
            .carryin(\PWMInstance0.un1_periodCounter_2_cry_11 ),
            .carryout(\PWMInstance0.un1_periodCounter_2_cry_12 ),
            .clk(N__38543),
            .ce(),
            .sr(N__35301));
    defparam \PWMInstance0.periodCounter_13_LC_7_17_5 .C_ON=1'b1;
    defparam \PWMInstance0.periodCounter_13_LC_7_17_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.periodCounter_13_LC_7_17_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance0.periodCounter_13_LC_7_17_5  (
            .in0(N__17288),
            .in1(N__18067),
            .in2(_gnd_net_),
            .in3(N__16074),
            .lcout(\PWMInstance0.periodCounterZ0Z_13 ),
            .ltout(),
            .carryin(\PWMInstance0.un1_periodCounter_2_cry_12 ),
            .carryout(\PWMInstance0.un1_periodCounter_2_cry_13 ),
            .clk(N__38543),
            .ce(),
            .sr(N__35301));
    defparam \PWMInstance0.periodCounter_14_LC_7_17_6 .C_ON=1'b1;
    defparam \PWMInstance0.periodCounter_14_LC_7_17_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.periodCounter_14_LC_7_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance0.periodCounter_14_LC_7_17_6  (
            .in0(_gnd_net_),
            .in1(N__17146),
            .in2(_gnd_net_),
            .in3(N__16071),
            .lcout(\PWMInstance0.periodCounterZ0Z_14 ),
            .ltout(),
            .carryin(\PWMInstance0.un1_periodCounter_2_cry_13 ),
            .carryout(\PWMInstance0.un1_periodCounter_2_cry_14 ),
            .clk(N__38543),
            .ce(),
            .sr(N__35301));
    defparam \PWMInstance0.periodCounter_15_LC_7_17_7 .C_ON=1'b1;
    defparam \PWMInstance0.periodCounter_15_LC_7_17_7 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.periodCounter_15_LC_7_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance0.periodCounter_15_LC_7_17_7  (
            .in0(_gnd_net_),
            .in1(N__17170),
            .in2(_gnd_net_),
            .in3(N__16068),
            .lcout(\PWMInstance0.periodCounterZ0Z_15 ),
            .ltout(),
            .carryin(\PWMInstance0.un1_periodCounter_2_cry_14 ),
            .carryout(\PWMInstance0.un1_periodCounter_2_cry_15 ),
            .clk(N__38543),
            .ce(),
            .sr(N__35301));
    defparam \PWMInstance0.periodCounter_16_LC_7_18_0 .C_ON=1'b0;
    defparam \PWMInstance0.periodCounter_16_LC_7_18_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.periodCounter_16_LC_7_18_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance0.periodCounter_16_LC_7_18_0  (
            .in0(N__17290),
            .in1(N__16060),
            .in2(_gnd_net_),
            .in3(N__16065),
            .lcout(\PWMInstance0.periodCounterZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38541),
            .ce(),
            .sr(N__35299));
    defparam \PWMInstance1.periodCounter_0_LC_8_1_0 .C_ON=1'b1;
    defparam \PWMInstance1.periodCounter_0_LC_8_1_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.periodCounter_0_LC_8_1_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance1.periodCounter_0_LC_8_1_0  (
            .in0(_gnd_net_),
            .in1(N__16042),
            .in2(N__16596),
            .in3(N__16595),
            .lcout(\PWMInstance1.periodCounterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_1_0_),
            .carryout(\PWMInstance1.un1_periodCounter_2_cry_0 ),
            .clk(N__38678),
            .ce(),
            .sr(N__35316));
    defparam \PWMInstance1.periodCounter_1_LC_8_1_1 .C_ON=1'b1;
    defparam \PWMInstance1.periodCounter_1_LC_8_1_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.periodCounter_1_LC_8_1_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance1.periodCounter_1_LC_8_1_1  (
            .in0(_gnd_net_),
            .in1(N__16618),
            .in2(_gnd_net_),
            .in3(N__16026),
            .lcout(\PWMInstance1.periodCounterZ0Z_1 ),
            .ltout(),
            .carryin(\PWMInstance1.un1_periodCounter_2_cry_0 ),
            .carryout(\PWMInstance1.un1_periodCounter_2_cry_1 ),
            .clk(N__38678),
            .ce(),
            .sr(N__35316));
    defparam \PWMInstance1.periodCounter_2_LC_8_1_2 .C_ON=1'b1;
    defparam \PWMInstance1.periodCounter_2_LC_8_1_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.periodCounter_2_LC_8_1_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance1.periodCounter_2_LC_8_1_2  (
            .in0(_gnd_net_),
            .in1(N__16023),
            .in2(_gnd_net_),
            .in3(N__16008),
            .lcout(\PWMInstance1.periodCounterZ0Z_2 ),
            .ltout(),
            .carryin(\PWMInstance1.un1_periodCounter_2_cry_1 ),
            .carryout(\PWMInstance1.un1_periodCounter_2_cry_2 ),
            .clk(N__38678),
            .ce(),
            .sr(N__35316));
    defparam \PWMInstance1.periodCounter_3_LC_8_1_3 .C_ON=1'b1;
    defparam \PWMInstance1.periodCounter_3_LC_8_1_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.periodCounter_3_LC_8_1_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance1.periodCounter_3_LC_8_1_3  (
            .in0(_gnd_net_),
            .in1(N__16241),
            .in2(_gnd_net_),
            .in3(N__16224),
            .lcout(\PWMInstance1.periodCounterZ0Z_3 ),
            .ltout(),
            .carryin(\PWMInstance1.un1_periodCounter_2_cry_2 ),
            .carryout(\PWMInstance1.un1_periodCounter_2_cry_3 ),
            .clk(N__38678),
            .ce(),
            .sr(N__35316));
    defparam \PWMInstance1.periodCounter_4_LC_8_1_4 .C_ON=1'b1;
    defparam \PWMInstance1.periodCounter_4_LC_8_1_4 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.periodCounter_4_LC_8_1_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance1.periodCounter_4_LC_8_1_4  (
            .in0(_gnd_net_),
            .in1(N__16221),
            .in2(_gnd_net_),
            .in3(N__16206),
            .lcout(\PWMInstance1.periodCounterZ0Z_4 ),
            .ltout(),
            .carryin(\PWMInstance1.un1_periodCounter_2_cry_3 ),
            .carryout(\PWMInstance1.un1_periodCounter_2_cry_4 ),
            .clk(N__38678),
            .ce(),
            .sr(N__35316));
    defparam \PWMInstance1.periodCounter_5_LC_8_1_5 .C_ON=1'b1;
    defparam \PWMInstance1.periodCounter_5_LC_8_1_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.periodCounter_5_LC_8_1_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance1.periodCounter_5_LC_8_1_5  (
            .in0(_gnd_net_),
            .in1(N__16202),
            .in2(_gnd_net_),
            .in3(N__16185),
            .lcout(\PWMInstance1.periodCounterZ0Z_5 ),
            .ltout(),
            .carryin(\PWMInstance1.un1_periodCounter_2_cry_4 ),
            .carryout(\PWMInstance1.un1_periodCounter_2_cry_5 ),
            .clk(N__38678),
            .ce(),
            .sr(N__35316));
    defparam \PWMInstance1.periodCounter_6_LC_8_1_6 .C_ON=1'b1;
    defparam \PWMInstance1.periodCounter_6_LC_8_1_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.periodCounter_6_LC_8_1_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance1.periodCounter_6_LC_8_1_6  (
            .in0(_gnd_net_),
            .in1(N__16172),
            .in2(_gnd_net_),
            .in3(N__16158),
            .lcout(\PWMInstance1.periodCounterZ0Z_6 ),
            .ltout(),
            .carryin(\PWMInstance1.un1_periodCounter_2_cry_5 ),
            .carryout(\PWMInstance1.un1_periodCounter_2_cry_6 ),
            .clk(N__38678),
            .ce(),
            .sr(N__35316));
    defparam \PWMInstance1.periodCounter_7_LC_8_1_7 .C_ON=1'b1;
    defparam \PWMInstance1.periodCounter_7_LC_8_1_7 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.periodCounter_7_LC_8_1_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance1.periodCounter_7_LC_8_1_7  (
            .in0(N__17000),
            .in1(N__16678),
            .in2(_gnd_net_),
            .in3(N__16155),
            .lcout(\PWMInstance1.periodCounterZ0Z_7 ),
            .ltout(),
            .carryin(\PWMInstance1.un1_periodCounter_2_cry_6 ),
            .carryout(\PWMInstance1.un1_periodCounter_2_cry_7 ),
            .clk(N__38678),
            .ce(),
            .sr(N__35316));
    defparam \PWMInstance1.periodCounter_8_LC_8_2_0 .C_ON=1'b1;
    defparam \PWMInstance1.periodCounter_8_LC_8_2_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.periodCounter_8_LC_8_2_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance1.periodCounter_8_LC_8_2_0  (
            .in0(_gnd_net_),
            .in1(N__16152),
            .in2(_gnd_net_),
            .in3(N__16134),
            .lcout(\PWMInstance1.periodCounterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_2_0_),
            .carryout(\PWMInstance1.un1_periodCounter_2_cry_8 ),
            .clk(N__38671),
            .ce(),
            .sr(N__35315));
    defparam \PWMInstance1.periodCounter_9_LC_8_2_1 .C_ON=1'b1;
    defparam \PWMInstance1.periodCounter_9_LC_8_2_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.periodCounter_9_LC_8_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance1.periodCounter_9_LC_8_2_1  (
            .in0(_gnd_net_),
            .in1(N__16130),
            .in2(_gnd_net_),
            .in3(N__16110),
            .lcout(\PWMInstance1.periodCounterZ0Z_9 ),
            .ltout(),
            .carryin(\PWMInstance1.un1_periodCounter_2_cry_8 ),
            .carryout(\PWMInstance1.un1_periodCounter_2_cry_9 ),
            .clk(N__38671),
            .ce(),
            .sr(N__35315));
    defparam \PWMInstance1.periodCounter_10_LC_8_2_2 .C_ON=1'b1;
    defparam \PWMInstance1.periodCounter_10_LC_8_2_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.periodCounter_10_LC_8_2_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance1.periodCounter_10_LC_8_2_2  (
            .in0(_gnd_net_),
            .in1(N__16103),
            .in2(_gnd_net_),
            .in3(N__16083),
            .lcout(\PWMInstance1.periodCounterZ0Z_10 ),
            .ltout(),
            .carryin(\PWMInstance1.un1_periodCounter_2_cry_9 ),
            .carryout(\PWMInstance1.un1_periodCounter_2_cry_10 ),
            .clk(N__38671),
            .ce(),
            .sr(N__35315));
    defparam \PWMInstance1.periodCounter_11_LC_8_2_3 .C_ON=1'b1;
    defparam \PWMInstance1.periodCounter_11_LC_8_2_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.periodCounter_11_LC_8_2_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance1.periodCounter_11_LC_8_2_3  (
            .in0(N__17002),
            .in1(N__16348),
            .in2(_gnd_net_),
            .in3(N__16326),
            .lcout(\PWMInstance1.periodCounterZ0Z_11 ),
            .ltout(),
            .carryin(\PWMInstance1.un1_periodCounter_2_cry_10 ),
            .carryout(\PWMInstance1.un1_periodCounter_2_cry_11 ),
            .clk(N__38671),
            .ce(),
            .sr(N__35315));
    defparam \PWMInstance1.periodCounter_12_LC_8_2_4 .C_ON=1'b1;
    defparam \PWMInstance1.periodCounter_12_LC_8_2_4 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.periodCounter_12_LC_8_2_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance1.periodCounter_12_LC_8_2_4  (
            .in0(N__17004),
            .in1(N__16322),
            .in2(_gnd_net_),
            .in3(N__16302),
            .lcout(\PWMInstance1.periodCounterZ0Z_12 ),
            .ltout(),
            .carryin(\PWMInstance1.un1_periodCounter_2_cry_11 ),
            .carryout(\PWMInstance1.un1_periodCounter_2_cry_12 ),
            .clk(N__38671),
            .ce(),
            .sr(N__35315));
    defparam \PWMInstance1.periodCounter_13_LC_8_2_5 .C_ON=1'b1;
    defparam \PWMInstance1.periodCounter_13_LC_8_2_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.periodCounter_13_LC_8_2_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance1.periodCounter_13_LC_8_2_5  (
            .in0(N__17003),
            .in1(N__16294),
            .in2(_gnd_net_),
            .in3(N__16275),
            .lcout(\PWMInstance1.periodCounterZ0Z_13 ),
            .ltout(),
            .carryin(\PWMInstance1.un1_periodCounter_2_cry_12 ),
            .carryout(\PWMInstance1.un1_periodCounter_2_cry_13 ),
            .clk(N__38671),
            .ce(),
            .sr(N__35315));
    defparam \PWMInstance1.periodCounter_14_LC_8_2_6 .C_ON=1'b1;
    defparam \PWMInstance1.periodCounter_14_LC_8_2_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.periodCounter_14_LC_8_2_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance1.periodCounter_14_LC_8_2_6  (
            .in0(_gnd_net_),
            .in1(N__16271),
            .in2(_gnd_net_),
            .in3(N__16251),
            .lcout(\PWMInstance1.periodCounterZ0Z_14 ),
            .ltout(),
            .carryin(\PWMInstance1.un1_periodCounter_2_cry_13 ),
            .carryout(\PWMInstance1.un1_periodCounter_2_cry_14 ),
            .clk(N__38671),
            .ce(),
            .sr(N__35315));
    defparam \PWMInstance1.periodCounter_15_LC_8_2_7 .C_ON=1'b1;
    defparam \PWMInstance1.periodCounter_15_LC_8_2_7 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.periodCounter_15_LC_8_2_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance1.periodCounter_15_LC_8_2_7  (
            .in0(_gnd_net_),
            .in1(N__16648),
            .in2(_gnd_net_),
            .in3(N__16248),
            .lcout(\PWMInstance1.periodCounterZ0Z_15 ),
            .ltout(),
            .carryin(\PWMInstance1.un1_periodCounter_2_cry_14 ),
            .carryout(\PWMInstance1.un1_periodCounter_2_cry_15 ),
            .clk(N__38671),
            .ce(),
            .sr(N__35315));
    defparam \PWMInstance1.periodCounter_16_LC_8_3_0 .C_ON=1'b0;
    defparam \PWMInstance1.periodCounter_16_LC_8_3_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.periodCounter_16_LC_8_3_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance1.periodCounter_16_LC_8_3_0  (
            .in0(N__17001),
            .in1(N__16702),
            .in2(_gnd_net_),
            .in3(N__16245),
            .lcout(\PWMInstance1.periodCounterZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38659),
            .ce(),
            .sr(N__35313));
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_1_c_LC_8_4_0 .C_ON=1'b1;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_1_c_LC_8_4_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_1_c_LC_8_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance5.un1_PWMPulseWidthCount_0_I_1_c_LC_8_4_0  (
            .in0(_gnd_net_),
            .in1(N__17907),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_4_0_),
            .carryout(\PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_9_c_LC_8_4_1 .C_ON=1'b1;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_9_c_LC_8_4_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_9_c_LC_8_4_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance5.un1_PWMPulseWidthCount_0_I_9_c_LC_8_4_1  (
            .in0(_gnd_net_),
            .in1(N__16962),
            .in2(N__32592),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_0 ),
            .carryout(\PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_15_c_LC_8_4_2 .C_ON=1'b1;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_15_c_LC_8_4_2 .SEQ_MODE=4'b0000;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_15_c_LC_8_4_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance5.un1_PWMPulseWidthCount_0_I_15_c_LC_8_4_2  (
            .in0(_gnd_net_),
            .in1(N__19272),
            .in2(N__32586),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_1 ),
            .carryout(\PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_27_c_LC_8_4_3 .C_ON=1'b1;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_27_c_LC_8_4_3 .SEQ_MODE=4'b0000;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_27_c_LC_8_4_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance5.un1_PWMPulseWidthCount_0_I_27_c_LC_8_4_3  (
            .in0(_gnd_net_),
            .in1(N__17883),
            .in2(N__32590),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_2 ),
            .carryout(\PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_45_c_LC_8_4_4 .C_ON=1'b1;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_45_c_LC_8_4_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_45_c_LC_8_4_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance5.un1_PWMPulseWidthCount_0_I_45_c_LC_8_4_4  (
            .in0(_gnd_net_),
            .in1(N__16416),
            .in2(N__32588),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_3 ),
            .carryout(\PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_33_c_LC_8_4_5 .C_ON=1'b1;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_33_c_LC_8_4_5 .SEQ_MODE=4'b0000;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_33_c_LC_8_4_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance5.un1_PWMPulseWidthCount_0_I_33_c_LC_8_4_5  (
            .in0(_gnd_net_),
            .in1(N__19143),
            .in2(N__32591),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_4 ),
            .carryout(\PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_39_c_LC_8_4_6 .C_ON=1'b1;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_39_c_LC_8_4_6 .SEQ_MODE=4'b0000;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_39_c_LC_8_4_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance5.un1_PWMPulseWidthCount_0_I_39_c_LC_8_4_6  (
            .in0(_gnd_net_),
            .in1(N__17220),
            .in2(N__32587),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_5 ),
            .carryout(\PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_21_c_LC_8_4_7 .C_ON=1'b1;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_21_c_LC_8_4_7 .SEQ_MODE=4'b0000;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_21_c_LC_8_4_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance5.un1_PWMPulseWidthCount_0_I_21_c_LC_8_4_7  (
            .in0(_gnd_net_),
            .in1(N__16932),
            .in2(N__32589),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_6 ),
            .carryout(\PWMInstance5.un1_PWMPulseWidthCount_0_data_tmp_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.out_LC_8_5_0 .C_ON=1'b0;
    defparam \PWMInstance5.out_LC_8_5_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.out_LC_8_5_0 .LUT_INIT=16'b1111101011110010;
    LogicCell40 \PWMInstance5.out_LC_8_5_0  (
            .in0(N__16385),
            .in1(N__19122),
            .in2(N__19461),
            .in3(N__16404),
            .lcout(PWM5_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38639),
            .ce(),
            .sr(N__35682));
    defparam \PWMInstance1.PWMPulseWidthCount_esr_12_LC_8_6_1 .C_ON=1'b0;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_12_LC_8_6_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_12_LC_8_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance1.PWMPulseWidthCount_esr_12_LC_8_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28875),
            .lcout(\PWMInstance1.PWMPulseWidthCountZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38628),
            .ce(N__16803),
            .sr(N__35685));
    defparam \PWMInstance1.PWMPulseWidthCount_esr_10_LC_8_6_4 .C_ON=1'b0;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_10_LC_8_6_4 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_10_LC_8_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance1.PWMPulseWidthCount_esr_10_LC_8_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36168),
            .lcout(\PWMInstance1.PWMPulseWidthCountZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38628),
            .ce(N__16803),
            .sr(N__35685));
    defparam \QuadInstance2.Quad_9_LC_8_7_0 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_9_LC_8_7_0 .SEQ_MODE=4'b1000;
    defparam \QuadInstance2.Quad_9_LC_8_7_0 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \QuadInstance2.Quad_9_LC_8_7_0  (
            .in0(_gnd_net_),
            .in1(N__28577),
            .in2(N__16359),
            .in3(N__22142),
            .lcout(dataRead2_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38617),
            .ce(),
            .sr(N__35691));
    defparam \QuadInstance2.Quad_10_LC_8_7_1 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_10_LC_8_7_1 .SEQ_MODE=4'b1000;
    defparam \QuadInstance2.Quad_10_LC_8_7_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance2.Quad_10_LC_8_7_1  (
            .in0(N__22139),
            .in1(N__36160),
            .in2(_gnd_net_),
            .in3(N__16434),
            .lcout(dataRead2_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38617),
            .ce(),
            .sr(N__35691));
    defparam \QuadInstance7.Quad_11_LC_8_7_2 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_11_LC_8_7_2 .SEQ_MODE=4'b1000;
    defparam \QuadInstance7.Quad_11_LC_8_7_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \QuadInstance7.Quad_11_LC_8_7_2  (
            .in0(N__36011),
            .in1(_gnd_net_),
            .in2(N__26037),
            .in3(N__17727),
            .lcout(dataRead7_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38617),
            .ce(),
            .sr(N__35691));
    defparam \QuadInstance4.Quad_9_LC_8_7_3 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_9_LC_8_7_3 .SEQ_MODE=4'b1000;
    defparam \QuadInstance4.Quad_9_LC_8_7_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance4.Quad_9_LC_8_7_3  (
            .in0(N__28578),
            .in1(N__29662),
            .in2(_gnd_net_),
            .in3(N__25050),
            .lcout(dataRead4_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38617),
            .ce(),
            .sr(N__35691));
    defparam \QuadInstance2.Quad_14_LC_8_7_4 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_14_LC_8_7_4 .SEQ_MODE=4'b1000;
    defparam \QuadInstance2.Quad_14_LC_8_7_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance2.Quad_14_LC_8_7_4  (
            .in0(N__34403),
            .in1(N__22141),
            .in2(_gnd_net_),
            .in3(N__16428),
            .lcout(dataRead2_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38617),
            .ce(),
            .sr(N__35691));
    defparam \QuadInstance1.Quad_2_LC_8_7_5 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_2_LC_8_7_5 .SEQ_MODE=4'b1000;
    defparam \QuadInstance1.Quad_2_LC_8_7_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance1.Quad_2_LC_8_7_5  (
            .in0(N__31593),
            .in1(N__24086),
            .in2(_gnd_net_),
            .in3(N__21633),
            .lcout(dataRead1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38617),
            .ce(),
            .sr(N__35691));
    defparam \QuadInstance7.Quad_12_LC_8_7_6 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_12_LC_8_7_6 .SEQ_MODE=4'b1000;
    defparam \QuadInstance7.Quad_12_LC_8_7_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance7.Quad_12_LC_8_7_6  (
            .in0(N__26004),
            .in1(N__28866),
            .in2(_gnd_net_),
            .in3(N__17706),
            .lcout(dataRead7_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38617),
            .ce(),
            .sr(N__35691));
    defparam \QuadInstance2.Quad_12_LC_8_7_7 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_12_LC_8_7_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance2.Quad_12_LC_8_7_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \QuadInstance2.Quad_12_LC_8_7_7  (
            .in0(N__22140),
            .in1(_gnd_net_),
            .in2(N__28874),
            .in3(N__16422),
            .lcout(dataRead2_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38617),
            .ce(),
            .sr(N__35691));
    defparam quadWrite_2_LC_8_8_0.C_ON=1'b0;
    defparam quadWrite_2_LC_8_8_0.SEQ_MODE=4'b1000;
    defparam quadWrite_2_LC_8_8_0.LUT_INIT=16'b0010000000000000;
    LogicCell40 quadWrite_2_LC_8_8_0 (
            .in0(N__33225),
            .in1(N__33848),
            .in2(N__33450),
            .in3(N__33652),
            .lcout(quadWriteZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38607),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNIB8VV2_4_LC_8_8_1 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_RNIB8VV2_4_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNIB8VV2_4_LC_8_8_1 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance7.Quad_RNIB8VV2_4_LC_8_8_1  (
            .in0(N__21465),
            .in1(N__25920),
            .in2(N__21800),
            .in3(N__16512),
            .lcout(\QuadInstance7.Quad_RNIB8VV2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam quadWrite_7_LC_8_8_2.C_ON=1'b0;
    defparam quadWrite_7_LC_8_8_2.SEQ_MODE=4'b1000;
    defparam quadWrite_7_LC_8_8_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 quadWrite_7_LC_8_8_2 (
            .in0(N__33847),
            .in1(N__33651),
            .in2(N__33451),
            .in3(N__23458),
            .lcout(quadWriteZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38607),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNIA7VV2_3_LC_8_8_3 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_RNIA7VV2_3_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNIA7VV2_3_LC_8_8_3 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance7.Quad_RNIA7VV2_3_LC_8_8_3  (
            .in0(N__27842),
            .in1(N__25919),
            .in2(N__21799),
            .in3(N__16510),
            .lcout(\QuadInstance7.Quad_RNIA7VV2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNIDAVV2_6_LC_8_8_4 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_RNIDAVV2_6_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNIDAVV2_6_LC_8_8_4 .LUT_INIT=16'b1111010100000000;
    LogicCell40 \QuadInstance7.Quad_RNIDAVV2_6_LC_8_8_4  (
            .in0(N__16513),
            .in1(N__27704),
            .in2(N__25971),
            .in3(N__21781),
            .lcout(\QuadInstance7.Quad_RNIDAVV2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNIEBVV2_7_LC_8_8_5 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_RNIEBVV2_7_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNIEBVV2_7_LC_8_8_5 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance7.Quad_RNIEBVV2_7_LC_8_8_5  (
            .in0(N__26271),
            .in1(N__25927),
            .in2(N__21801),
            .in3(N__16514),
            .lcout(\QuadInstance7.Quad_RNIEBVV2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNIC9VV2_5_LC_8_8_6 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_RNIC9VV2_5_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNIC9VV2_5_LC_8_8_6 .LUT_INIT=16'b1111010100000000;
    LogicCell40 \QuadInstance7.Quad_RNIC9VV2_5_LC_8_8_6  (
            .in0(N__16511),
            .in1(N__36746),
            .in2(N__25970),
            .in3(N__21777),
            .lcout(\QuadInstance7.Quad_RNIC9VV2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNIOIKU2_10_LC_8_9_0 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_RNIOIKU2_10_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNIOIKU2_10_LC_8_9_0 .LUT_INIT=16'b1100000011001100;
    LogicCell40 \QuadInstance7.Quad_RNIOIKU2_10_LC_8_9_0  (
            .in0(N__34650),
            .in1(N__21787),
            .in2(N__25973),
            .in3(N__16508),
            .lcout(\QuadInstance7.Quad_RNIOIKU2Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.delayedCh_B_RNI2N241_2_LC_8_9_1 .C_ON=1'b0;
    defparam \QuadInstance7.delayedCh_B_RNI2N241_2_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.delayedCh_B_RNI2N241_2_LC_8_9_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \QuadInstance7.delayedCh_B_RNI2N241_2_LC_8_9_1  (
            .in0(N__34470),
            .in1(N__16841),
            .in2(_gnd_net_),
            .in3(N__16462),
            .lcout(\QuadInstance7.un1_count_enable_i_a2_0_1 ),
            .ltout(\QuadInstance7.un1_count_enable_i_a2_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNI96VV2_2_LC_8_9_2 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_RNI96VV2_2_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNI96VV2_2_LC_8_9_2 .LUT_INIT=16'b1100111100000000;
    LogicCell40 \QuadInstance7.Quad_RNI96VV2_2_LC_8_9_2  (
            .in0(N__30386),
            .in1(N__25918),
            .in2(N__16440),
            .in3(N__21782),
            .lcout(\QuadInstance7.Quad_RNI96VV2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.delayedCh_A_RNI8MRP1_2_LC_8_9_3 .C_ON=1'b0;
    defparam \QuadInstance7.delayedCh_A_RNI8MRP1_2_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.delayedCh_A_RNI8MRP1_2_LC_8_9_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \QuadInstance7.delayedCh_A_RNI8MRP1_2_LC_8_9_3  (
            .in0(N__16853),
            .in1(N__16463),
            .in2(N__16449),
            .in3(N__16842),
            .lcout(\QuadInstance7.count_enable ),
            .ltout(\QuadInstance7.count_enable_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNI85VV2_1_LC_8_9_4 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_RNI85VV2_1_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNI85VV2_1_LC_8_9_4 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance7.Quad_RNI85VV2_1_LC_8_9_4  (
            .in0(N__25841),
            .in1(N__25917),
            .in2(N__16437),
            .in3(N__16505),
            .lcout(\QuadInstance7.Quad_RNI85VV2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNIFCVV2_8_LC_8_9_5 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_RNIFCVV2_8_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNIFCVV2_8_LC_8_9_5 .LUT_INIT=16'b1101000011010000;
    LogicCell40 \QuadInstance7.Quad_RNIFCVV2_8_LC_8_9_5  (
            .in0(N__16506),
            .in1(N__25928),
            .in2(N__21802),
            .in3(N__37613),
            .lcout(\QuadInstance7.Quad_RNIFCVV2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNIGDVV2_9_LC_8_9_6 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_RNIGDVV2_9_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNIGDVV2_9_LC_8_9_6 .LUT_INIT=16'b1100000011001100;
    LogicCell40 \QuadInstance7.Quad_RNIGDVV2_9_LC_8_9_6  (
            .in0(N__25392),
            .in1(N__21786),
            .in2(N__25972),
            .in3(N__16507),
            .lcout(\QuadInstance7.Quad_RNIGDVV2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNIRLKU2_13_LC_8_9_7 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_RNIRLKU2_13_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNIRLKU2_13_LC_8_9_7 .LUT_INIT=16'b1101000011010000;
    LogicCell40 \QuadInstance7.Quad_RNIRLKU2_13_LC_8_9_7  (
            .in0(N__16509),
            .in1(N__25935),
            .in2(N__21803),
            .in3(N__26112),
            .lcout(\QuadInstance7.Quad_RNIRLKU2Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNISMKU2_14_LC_8_10_0 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_RNISMKU2_14_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNISMKU2_14_LC_8_10_0 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \QuadInstance7.Quad_RNISMKU2_14_LC_8_10_0  (
            .in0(N__16521),
            .in1(N__25976),
            .in2(N__20283),
            .in3(N__21794),
            .lcout(\QuadInstance7.Quad_RNISMKU2Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.delayedCh_B_1_LC_8_10_1 .C_ON=1'b0;
    defparam \QuadInstance7.delayedCh_B_1_LC_8_10_1 .SEQ_MODE=4'b1000;
    defparam \QuadInstance7.delayedCh_B_1_LC_8_10_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \QuadInstance7.delayedCh_B_1_LC_8_10_1  (
            .in0(N__17418),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\QuadInstance7.delayedCh_BZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38587),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNIPJKU2_11_LC_8_10_2 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_RNIPJKU2_11_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNIPJKU2_11_LC_8_10_2 .LUT_INIT=16'b1100111100000000;
    LogicCell40 \QuadInstance7.Quad_RNIPJKU2_11_LC_8_10_2  (
            .in0(N__20877),
            .in1(N__25974),
            .in2(N__16523),
            .in3(N__21792),
            .lcout(\QuadInstance7.Quad_RNIPJKU2Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.delayedCh_A_1_LC_8_10_3 .C_ON=1'b0;
    defparam \QuadInstance7.delayedCh_A_1_LC_8_10_3 .SEQ_MODE=4'b1000;
    defparam \QuadInstance7.delayedCh_A_1_LC_8_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance7.delayedCh_A_1_LC_8_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29694),
            .lcout(\QuadInstance7.delayedCh_AZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38587),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNIQKKU2_12_LC_8_10_4 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_RNIQKKU2_12_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNIQKKU2_12_LC_8_10_4 .LUT_INIT=16'b1100111100000000;
    LogicCell40 \QuadInstance7.Quad_RNIQKKU2_12_LC_8_10_4  (
            .in0(N__22262),
            .in1(N__25975),
            .in2(N__16524),
            .in3(N__21793),
            .lcout(\QuadInstance7.Quad_RNIQKKU2Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwmWrite_1_LC_8_10_5.C_ON=1'b0;
    defparam pwmWrite_1_LC_8_10_5.SEQ_MODE=4'b1000;
    defparam pwmWrite_1_LC_8_10_5.LUT_INIT=16'b0000000000000010;
    LogicCell40 pwmWrite_1_LC_8_10_5 (
            .in0(N__23451),
            .in1(N__33830),
            .in2(N__33442),
            .in3(N__33666),
            .lcout(pwmWriteZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38587),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.delayedCh_A_2_LC_8_10_6 .C_ON=1'b0;
    defparam \QuadInstance7.delayedCh_A_2_LC_8_10_6 .SEQ_MODE=4'b1000;
    defparam \QuadInstance7.delayedCh_A_2_LC_8_10_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \QuadInstance7.delayedCh_A_2_LC_8_10_6  (
            .in0(N__16464),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\QuadInstance7.delayedCh_AZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38587),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.delayedCh_B_2_LC_8_10_7 .C_ON=1'b0;
    defparam \QuadInstance7.delayedCh_B_2_LC_8_10_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance7.delayedCh_B_2_LC_8_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance7.delayedCh_B_2_LC_8_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16854),
            .lcout(\QuadInstance7.delayedCh_BZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38587),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance1.out_RNO_0_LC_8_11_0 .C_ON=1'b0;
    defparam \PWMInstance1.out_RNO_0_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance1.out_RNO_0_LC_8_11_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \PWMInstance1.out_RNO_0_LC_8_11_0  (
            .in0(N__17823),
            .in1(N__16735),
            .in2(N__16707),
            .in3(N__16720),
            .lcout(\PWMInstance1.un1_periodCounter12_1_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance1.clkCount_0_LC_8_11_1 .C_ON=1'b0;
    defparam \PWMInstance1.clkCount_0_LC_8_11_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.clkCount_0_LC_8_11_1 .LUT_INIT=16'b1010101000000101;
    LogicCell40 \PWMInstance1.clkCount_0_LC_8_11_1  (
            .in0(N__16721),
            .in1(_gnd_net_),
            .in2(N__16742),
            .in3(N__16754),
            .lcout(\PWMInstance1.clkCountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38576),
            .ce(),
            .sr(N__35720));
    defparam \PWMInstance1.PWMPulseWidthCount_esr_ctle_15_LC_8_11_2 .C_ON=1'b0;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_ctle_15_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \PWMInstance1.PWMPulseWidthCount_esr_ctle_15_LC_8_11_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \PWMInstance1.PWMPulseWidthCount_esr_ctle_15_LC_8_11_2  (
            .in0(N__16753),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35825),
            .lcout(\PWMInstance1.pwmWrite_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance1.clkCount_1_LC_8_11_3 .C_ON=1'b0;
    defparam \PWMInstance1.clkCount_1_LC_8_11_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance1.clkCount_1_LC_8_11_3 .LUT_INIT=16'b1111000000001010;
    LogicCell40 \PWMInstance1.clkCount_1_LC_8_11_3  (
            .in0(N__16722),
            .in1(_gnd_net_),
            .in2(N__16743),
            .in3(N__16755),
            .lcout(\PWMInstance1.clkCountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38576),
            .ce(),
            .sr(N__35720));
    defparam \PWMInstance1.clkCount_RNISE5O_0_LC_8_11_4 .C_ON=1'b0;
    defparam \PWMInstance1.clkCount_RNISE5O_0_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance1.clkCount_RNISE5O_0_LC_8_11_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \PWMInstance1.clkCount_RNISE5O_0_LC_8_11_4  (
            .in0(N__17822),
            .in1(N__16734),
            .in2(_gnd_net_),
            .in3(N__16719),
            .lcout(\PWMInstance1.periodCounter12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance1.periodCounter_RNI4EVP_16_LC_8_11_5 .C_ON=1'b0;
    defparam \PWMInstance1.periodCounter_RNI4EVP_16_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \PWMInstance1.periodCounter_RNI4EVP_16_LC_8_11_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \PWMInstance1.periodCounter_RNI4EVP_16_LC_8_11_5  (
            .in0(_gnd_net_),
            .in1(N__16703),
            .in2(_gnd_net_),
            .in3(N__16686),
            .lcout(),
            .ltout(\PWMInstance1.un1_periodCounter12_1_0_a2_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance1.periodCounter_RNIT34C2_1_LC_8_11_6 .C_ON=1'b0;
    defparam \PWMInstance1.periodCounter_RNIT34C2_1_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \PWMInstance1.periodCounter_RNIT34C2_1_LC_8_11_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \PWMInstance1.periodCounter_RNIT34C2_1_LC_8_11_6  (
            .in0(N__16655),
            .in1(N__16626),
            .in2(N__16599),
            .in3(N__16580),
            .lcout(),
            .ltout(\PWMInstance1.un1_periodCounter12_1_0_a2_0_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance1.periodCounter_RNIOA6I7_0_LC_8_11_7 .C_ON=1'b0;
    defparam \PWMInstance1.periodCounter_RNIOA6I7_0_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \PWMInstance1.periodCounter_RNIOA6I7_0_LC_8_11_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \PWMInstance1.periodCounter_RNIOA6I7_0_LC_8_11_7  (
            .in0(N__16569),
            .in1(N__16554),
            .in2(N__16542),
            .in3(N__16539),
            .lcout(\PWMInstance1.out_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_8_12_1 .C_ON=1'b0;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_8_12_1 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance5.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_8_12_1  (
            .in0(N__16947),
            .in1(N__16953),
            .in2(N__19346),
            .in3(N__19256),
            .lcout(\PWMInstance5.un1_PWMPulseWidthCount_0_I_9_c_RNO_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.PWMPulseWidthCount_esr_2_LC_8_12_2 .C_ON=1'b0;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_2_LC_8_12_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_2_LC_8_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance5.PWMPulseWidthCount_esr_2_LC_8_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31591),
            .lcout(\PWMInstance5.PWMPulseWidthCountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38566),
            .ce(N__19635),
            .sr(N__35728));
    defparam \PWMInstance5.PWMPulseWidthCount_esr_3_LC_8_12_3 .C_ON=1'b0;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_3_LC_8_12_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_3_LC_8_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance5.PWMPulseWidthCount_esr_3_LC_8_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32085),
            .lcout(\PWMInstance5.PWMPulseWidthCountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38566),
            .ce(N__19635),
            .sr(N__35728));
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_8_12_4 .C_ON=1'b0;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_8_12_4 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \PWMInstance5.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_8_12_4  (
            .in0(N__16941),
            .in1(N__16920),
            .in2(N__19524),
            .in3(N__19238),
            .lcout(\PWMInstance5.un1_PWMPulseWidthCount_0_I_21_c_RNO_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.PWMPulseWidthCount_esr_15_LC_8_12_6 .C_ON=1'b0;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_15_LC_8_12_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_15_LC_8_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance5.PWMPulseWidthCount_esr_15_LC_8_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31871),
            .lcout(\PWMInstance5.PWMPulseWidthCountZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38566),
            .ce(N__19635),
            .sr(N__35728));
    defparam pwmWrite_0_LC_8_13_0.C_ON=1'b0;
    defparam pwmWrite_0_LC_8_13_0.SEQ_MODE=4'b1000;
    defparam pwmWrite_0_LC_8_13_0.LUT_INIT=16'b0000000100000000;
    LogicCell40 pwmWrite_0_LC_8_13_0 (
            .in0(N__33849),
            .in1(N__33672),
            .in2(N__33452),
            .in3(N__33224),
            .lcout(pwmWriteZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38560),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_8_13_1 .C_ON=1'b0;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_8_13_1 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \PWMInstance0.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_8_13_1  (
            .in0(N__18140),
            .in1(N__16914),
            .in2(N__16908),
            .in3(N__16881),
            .lcout(\PWMInstance0.un1_PWMPulseWidthCount_0_I_45_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance0.PWMPulseWidthCount_esr_ctle_15_LC_8_13_3 .C_ON=1'b0;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_ctle_15_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_ctle_15_LC_8_13_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \PWMInstance0.PWMPulseWidthCount_esr_ctle_15_LC_8_13_3  (
            .in0(N__35826),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16865),
            .lcout(\PWMInstance0.pwmWrite_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_8_13_4 .C_ON=1'b0;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_8_13_4 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance5.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_8_13_4  (
            .in0(N__18210),
            .in1(N__17232),
            .in2(N__18177),
            .in3(N__19220),
            .lcout(\PWMInstance5.un1_PWMPulseWidthCount_0_I_39_c_RNO_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_8_13_7 .C_ON=1'b0;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_8_13_7 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \PWMInstance0.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_8_13_7  (
            .in0(N__18261),
            .in1(N__17208),
            .in2(N__18111),
            .in3(N__17202),
            .lcout(\PWMInstance0.un1_PWMPulseWidthCount_0_I_27_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_8_14_0 .C_ON=1'b0;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_8_14_0 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance0.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_8_14_0  (
            .in0(N__17118),
            .in1(N__17124),
            .in2(N__17178),
            .in3(N__17151),
            .lcout(\PWMInstance0.un1_PWMPulseWidthCount_0_I_21_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance0.PWMPulseWidthCount_esr_14_LC_8_14_1 .C_ON=1'b0;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_14_LC_8_14_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_14_LC_8_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance0.PWMPulseWidthCount_esr_14_LC_8_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34378),
            .lcout(\PWMInstance0.PWMPulseWidthCountZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38553),
            .ce(N__18234),
            .sr(N__35743));
    defparam \PWMInstance0.PWMPulseWidthCount_esr_15_LC_8_14_2 .C_ON=1'b0;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_15_LC_8_14_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_15_LC_8_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance0.PWMPulseWidthCount_esr_15_LC_8_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31878),
            .lcout(\PWMInstance0.PWMPulseWidthCountZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38553),
            .ce(N__18234),
            .sr(N__35743));
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_8_14_3 .C_ON=1'b0;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_8_14_3 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \PWMInstance0.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_8_14_3  (
            .in0(N__17111),
            .in1(N__17046),
            .in2(N__17087),
            .in3(N__17058),
            .lcout(\PWMInstance0.un1_PWMPulseWidthCount_0_I_33_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance0.PWMPulseWidthCount_esr_11_LC_8_14_5 .C_ON=1'b0;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_11_LC_8_14_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_11_LC_8_14_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \PWMInstance0.PWMPulseWidthCount_esr_11_LC_8_14_5  (
            .in0(_gnd_net_),
            .in1(N__35998),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PWMInstance0.PWMPulseWidthCountZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38553),
            .ce(N__18234),
            .sr(N__35743));
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_8_14_6 .C_ON=1'b0;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_8_14_6 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance0.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_8_14_6  (
            .in0(N__17040),
            .in1(N__17034),
            .in2(N__18077),
            .in3(N__17028),
            .lcout(\PWMInstance0.un1_PWMPulseWidthCount_0_I_39_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_1_c_LC_8_15_0 .C_ON=1'b1;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_1_c_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_1_c_LC_8_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance0.un1_PWMPulseWidthCount_0_I_1_c_LC_8_15_0  (
            .in0(_gnd_net_),
            .in1(N__17988),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_15_0_),
            .carryout(\PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_9_c_LC_8_15_1 .C_ON=1'b1;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_9_c_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_9_c_LC_8_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance0.un1_PWMPulseWidthCount_0_I_9_c_LC_8_15_1  (
            .in0(_gnd_net_),
            .in1(N__17346),
            .in2(N__32572),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_0 ),
            .carryout(\PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_15_c_LC_8_15_2 .C_ON=1'b1;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_15_c_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_15_c_LC_8_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance0.un1_PWMPulseWidthCount_0_I_15_c_LC_8_15_2  (
            .in0(_gnd_net_),
            .in1(N__17340),
            .in2(N__32566),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_1 ),
            .carryout(\PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_27_c_LC_8_15_3 .C_ON=1'b1;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_27_c_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_27_c_LC_8_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance0.un1_PWMPulseWidthCount_0_I_27_c_LC_8_15_3  (
            .in0(_gnd_net_),
            .in1(N__17334),
            .in2(N__32570),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_2 ),
            .carryout(\PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_45_c_LC_8_15_4 .C_ON=1'b1;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_45_c_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_45_c_LC_8_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance0.un1_PWMPulseWidthCount_0_I_45_c_LC_8_15_4  (
            .in0(_gnd_net_),
            .in1(N__17325),
            .in2(N__32568),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_3 ),
            .carryout(\PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_33_c_LC_8_15_5 .C_ON=1'b1;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_33_c_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_33_c_LC_8_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance0.un1_PWMPulseWidthCount_0_I_33_c_LC_8_15_5  (
            .in0(_gnd_net_),
            .in1(N__17316),
            .in2(N__32571),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_4 ),
            .carryout(\PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_39_c_LC_8_15_6 .C_ON=1'b1;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_39_c_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_39_c_LC_8_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance0.un1_PWMPulseWidthCount_0_I_39_c_LC_8_15_6  (
            .in0(_gnd_net_),
            .in1(N__17310),
            .in2(N__32567),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_5 ),
            .carryout(\PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_21_c_LC_8_15_7 .C_ON=1'b1;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_21_c_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_21_c_LC_8_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance0.un1_PWMPulseWidthCount_0_I_21_c_LC_8_15_7  (
            .in0(_gnd_net_),
            .in1(N__17304),
            .in2(N__32569),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_6 ),
            .carryout(\PWMInstance0.un1_PWMPulseWidthCount_0_data_tmp_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance0.out_LC_8_16_0 .C_ON=1'b0;
    defparam \PWMInstance0.out_LC_8_16_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.out_LC_8_16_0 .LUT_INIT=16'b1111101011110010;
    LogicCell40 \PWMInstance0.out_LC_8_16_0  (
            .in0(N__17243),
            .in1(N__17298),
            .in2(N__17292),
            .in3(N__17253),
            .lcout(PWM0_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38546),
            .ce(),
            .sr(N__35755));
    defparam \QuadInstance7.delayedCh_B_0_LC_8_19_0 .C_ON=1'b0;
    defparam \QuadInstance7.delayedCh_B_0_LC_8_19_0 .SEQ_MODE=4'b1000;
    defparam \QuadInstance7.delayedCh_B_0_LC_8_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance7.delayedCh_B_0_LC_8_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17436),
            .lcout(\QuadInstance7.delayedCh_BZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38542),
            .ce(),
            .sr(_gnd_net_));
    defparam PWM0_obufLegalizeSB_DFF_LC_8_20_0.C_ON=1'b0;
    defparam PWM0_obufLegalizeSB_DFF_LC_8_20_0.SEQ_MODE=4'b1000;
    defparam PWM0_obufLegalizeSB_DFF_LC_8_20_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 PWM0_obufLegalizeSB_DFF_LC_8_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PWM0_obufLegalizeSB_DFFNet),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36936),
            .ce(),
            .sr(_gnd_net_));
    defparam PWM1_obufLegalizeSB_DFF_LC_8_20_1.C_ON=1'b0;
    defparam PWM1_obufLegalizeSB_DFF_LC_8_20_1.SEQ_MODE=4'b1000;
    defparam PWM1_obufLegalizeSB_DFF_LC_8_20_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 PWM1_obufLegalizeSB_DFF_LC_8_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PWM1_obufLegalizeSB_DFFNet),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36936),
            .ce(),
            .sr(_gnd_net_));
    defparam PWM6_obufLegalizeSB_DFF_LC_8_20_2.C_ON=1'b0;
    defparam PWM6_obufLegalizeSB_DFF_LC_8_20_2.SEQ_MODE=4'b1000;
    defparam PWM6_obufLegalizeSB_DFF_LC_8_20_2.LUT_INIT=16'b1111111111111111;
    LogicCell40 PWM6_obufLegalizeSB_DFF_LC_8_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PWM6_obufLegalizeSB_DFFNet),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36936),
            .ce(),
            .sr(_gnd_net_));
    defparam PWM7_obufLegalizeSB_DFF_LC_8_20_3.C_ON=1'b0;
    defparam PWM7_obufLegalizeSB_DFF_LC_8_20_3.SEQ_MODE=4'b1000;
    defparam PWM7_obufLegalizeSB_DFF_LC_8_20_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 PWM7_obufLegalizeSB_DFF_LC_8_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PWM7_obufLegalizeSB_DFFNet),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36936),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.delayedCh_B_0_LC_9_2_4 .C_ON=1'b0;
    defparam \QuadInstance3.delayedCh_B_0_LC_9_2_4 .SEQ_MODE=4'b1000;
    defparam \QuadInstance3.delayedCh_B_0_LC_9_2_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \QuadInstance3.delayedCh_B_0_LC_9_2_4  (
            .in0(N__17385),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\QuadInstance3.delayedCh_BZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38679),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_4_LC_9_3_5 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_4_LC_9_3_5 .SEQ_MODE=4'b1000;
    defparam \QuadInstance2.Quad_4_LC_9_3_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance2.Quad_4_LC_9_3_5  (
            .in0(N__36521),
            .in1(N__22171),
            .in2(_gnd_net_),
            .in3(N__17376),
            .lcout(dataRead2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38672),
            .ce(),
            .sr(N__35681));
    defparam \QuadInstance5.delayedCh_A_1_LC_9_4_1 .C_ON=1'b0;
    defparam \QuadInstance5.delayedCh_A_1_LC_9_4_1 .SEQ_MODE=4'b1000;
    defparam \QuadInstance5.delayedCh_A_1_LC_9_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance5.delayedCh_A_1_LC_9_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17352),
            .lcout(\QuadInstance5.delayedCh_AZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38660),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.delayedCh_A_0_LC_9_4_4 .C_ON=1'b0;
    defparam \QuadInstance5.delayedCh_A_0_LC_9_4_4 .SEQ_MODE=4'b1000;
    defparam \QuadInstance5.delayedCh_A_0_LC_9_4_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance5.delayedCh_A_0_LC_9_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17364),
            .lcout(\QuadInstance5.delayedCh_AZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38660),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNI07LI2_9_LC_9_5_0 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_RNI07LI2_9_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNI07LI2_9_LC_9_5_0 .LUT_INIT=16'b1100111100000000;
    LogicCell40 \QuadInstance5.Quad_RNI07LI2_9_LC_9_5_0  (
            .in0(N__25514),
            .in1(N__25727),
            .in2(N__17500),
            .in3(N__18368),
            .lcout(\QuadInstance5.Quad_RNI07LI2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.delayedCh_B_RNIUQSQ_2_LC_9_5_1 .C_ON=1'b0;
    defparam \QuadInstance5.delayedCh_B_RNIUQSQ_2_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.delayedCh_B_RNIUQSQ_2_LC_9_5_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \QuadInstance5.delayedCh_B_RNIUQSQ_2_LC_9_5_1  (
            .in0(N__34500),
            .in1(N__18407),
            .in2(_gnd_net_),
            .in3(N__18433),
            .lcout(\QuadInstance5.un1_count_enable_i_a2_0_1 ),
            .ltout(\QuadInstance5.un1_count_enable_i_a2_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNIPVKI2_2_LC_9_5_2 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_RNIPVKI2_2_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNIPVKI2_2_LC_9_5_2 .LUT_INIT=16'b1100111100000000;
    LogicCell40 \QuadInstance5.Quad_RNIPVKI2_2_LC_9_5_2  (
            .in0(N__30530),
            .in1(N__25723),
            .in2(N__17439),
            .in3(N__18360),
            .lcout(\QuadInstance5.Quad_RNIPVKI2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNIQ0LI2_3_LC_9_5_4 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_RNIQ0LI2_3_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNIQ0LI2_3_LC_9_5_4 .LUT_INIT=16'b1100111100000000;
    LogicCell40 \QuadInstance5.Quad_RNIQ0LI2_3_LC_9_5_4  (
            .in0(N__27918),
            .in1(N__25724),
            .in2(N__17499),
            .in3(N__18364),
            .lcout(\QuadInstance5.Quad_RNIQ0LI2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNIR1LI2_4_LC_9_5_5 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_RNIR1LI2_4_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNIR1LI2_4_LC_9_5_5 .LUT_INIT=16'b1010000011110000;
    LogicCell40 \QuadInstance5.Quad_RNIR1LI2_4_LC_9_5_5  (
            .in0(N__25725),
            .in1(N__21326),
            .in2(N__18382),
            .in3(N__17478),
            .lcout(\QuadInstance5.Quad_RNIR1LI2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNIS2LI2_5_LC_9_5_7 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_RNIS2LI2_5_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNIS2LI2_5_LC_9_5_7 .LUT_INIT=16'b1010000011110000;
    LogicCell40 \QuadInstance5.Quad_RNIS2LI2_5_LC_9_5_7  (
            .in0(N__25726),
            .in1(N__36871),
            .in2(N__18383),
            .in3(N__17482),
            .lcout(\QuadInstance5.Quad_RNIS2LI2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNI8AQ82_10_LC_9_6_0 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_RNI8AQ82_10_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNI8AQ82_10_LC_9_6_0 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \QuadInstance5.Quad_RNI8AQ82_10_LC_9_6_0  (
            .in0(N__25722),
            .in1(N__17486),
            .in2(N__35024),
            .in3(N__18358),
            .lcout(\QuadInstance5.Quad_RNI8AQ82Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNI9BQ82_11_LC_9_6_1 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_RNI9BQ82_11_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNI9BQ82_11_LC_9_6_1 .LUT_INIT=16'b1000101010001010;
    LogicCell40 \QuadInstance5.Quad_RNI9BQ82_11_LC_9_6_1  (
            .in0(N__18359),
            .in1(N__25721),
            .in2(N__17501),
            .in3(N__20112),
            .lcout(\QuadInstance5.Quad_RNI9BQ82Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam quadWrite_5_LC_9_6_2.C_ON=1'b0;
    defparam quadWrite_5_LC_9_6_2.SEQ_MODE=4'b1000;
    defparam quadWrite_5_LC_9_6_2.LUT_INIT=16'b0010000000000000;
    LogicCell40 quadWrite_5_LC_9_6_2 (
            .in0(N__33827),
            .in1(N__33639),
            .in2(N__33466),
            .in3(N__23459),
            .lcout(quadWriteZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38640),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNIT3LI2_6_LC_9_6_3 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_RNIT3LI2_6_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNIT3LI2_6_LC_9_6_3 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance5.Quad_RNIT3LI2_6_LC_9_6_3  (
            .in0(N__25281),
            .in1(N__25716),
            .in2(N__18380),
            .in3(N__17476),
            .lcout(\QuadInstance5.Quad_RNIT3LI2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNIU4LI2_7_LC_9_6_4 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_RNIU4LI2_7_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNIU4LI2_7_LC_9_6_4 .LUT_INIT=16'b1111010100000000;
    LogicCell40 \QuadInstance5.Quad_RNIU4LI2_7_LC_9_6_4  (
            .in0(N__17475),
            .in1(N__25607),
            .in2(N__25757),
            .in3(N__18351),
            .lcout(\QuadInstance5.Quad_RNIU4LI2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNIV5LI2_8_LC_9_6_5 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_RNIV5LI2_8_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNIV5LI2_8_LC_9_6_5 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance5.Quad_RNIV5LI2_8_LC_9_6_5  (
            .in0(N__36984),
            .in1(N__25720),
            .in2(N__18381),
            .in3(N__17477),
            .lcout(\QuadInstance5.Quad_RNIV5LI2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_RNIJ03G2_13_LC_9_6_6 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_RNIJ03G2_13_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \QuadInstance2.Quad_RNIJ03G2_13_LC_9_6_6 .LUT_INIT=16'b1100111100000000;
    LogicCell40 \QuadInstance2.Quad_RNIJ03G2_13_LC_9_6_6  (
            .in0(N__19974),
            .in1(N__22143),
            .in2(N__17601),
            .in3(N__18530),
            .lcout(\QuadInstance2.Quad_RNIJ03G2Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNIOUKI2_1_LC_9_6_7 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_RNIOUKI2_1_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNIOUKI2_1_LC_9_6_7 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance5.Quad_RNIOUKI2_1_LC_9_6_7  (
            .in0(N__23858),
            .in1(N__25715),
            .in2(N__18379),
            .in3(N__17474),
            .lcout(\QuadInstance5.Quad_RNIOUKI2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNIACQ82_12_LC_9_7_0 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_RNIACQ82_12_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNIACQ82_12_LC_9_7_0 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \QuadInstance5.Quad_RNIACQ82_12_LC_9_7_0  (
            .in0(N__25728),
            .in1(N__17503),
            .in2(N__22385),
            .in3(N__18387),
            .lcout(\QuadInstance5.Quad_RNIACQ82Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNIBDQ82_13_LC_9_7_1 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_RNIBDQ82_13_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNIBDQ82_13_LC_9_7_1 .LUT_INIT=16'b1111000001010000;
    LogicCell40 \QuadInstance5.Quad_RNIBDQ82_13_LC_9_7_1  (
            .in0(N__17502),
            .in1(N__20008),
            .in2(N__18392),
            .in3(N__25729),
            .lcout(\QuadInstance5.Quad_RNIBDQ82Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNICEQ82_14_LC_9_7_2 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_RNICEQ82_14_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNICEQ82_14_LC_9_7_2 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \QuadInstance5.Quad_RNICEQ82_14_LC_9_7_2  (
            .in0(N__25730),
            .in1(N__18388),
            .in2(N__28222),
            .in3(N__17504),
            .lcout(\QuadInstance5.Quad_RNICEQ82Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNO_0_15_LC_9_7_3 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_RNO_0_15_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNO_0_15_LC_9_7_3 .LUT_INIT=16'b0011110010011100;
    LogicCell40 \QuadInstance5.Quad_RNO_0_15_LC_9_7_3  (
            .in0(N__17505),
            .in1(N__24242),
            .in2(N__18393),
            .in3(N__25731),
            .lcout(\QuadInstance5.un1_Quad_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_12_LC_9_7_4 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_12_LC_9_7_4 .SEQ_MODE=4'b1000;
    defparam \QuadInstance5.Quad_12_LC_9_7_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance5.Quad_12_LC_9_7_4  (
            .in0(N__25732),
            .in1(N__28847),
            .in2(_gnd_net_),
            .in3(N__18543),
            .lcout(dataRead5_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38629),
            .ce(),
            .sr(N__35698));
    defparam \QuadInstance5.Quad_13_LC_9_7_5 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_13_LC_9_7_5 .SEQ_MODE=4'b1000;
    defparam \QuadInstance5.Quad_13_LC_9_7_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance5.Quad_13_LC_9_7_5  (
            .in0(N__28719),
            .in1(N__25734),
            .in2(_gnd_net_),
            .in3(N__18705),
            .lcout(dataRead5_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38629),
            .ce(),
            .sr(N__35698));
    defparam \QuadInstance5.Quad_14_LC_9_7_6 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_14_LC_9_7_6 .SEQ_MODE=4'b1000;
    defparam \QuadInstance5.Quad_14_LC_9_7_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance5.Quad_14_LC_9_7_6  (
            .in0(N__25733),
            .in1(N__34402),
            .in2(_gnd_net_),
            .in3(N__18690),
            .lcout(dataRead5_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38629),
            .ce(),
            .sr(N__35698));
    defparam \QuadInstance5.Quad_1_LC_9_7_7 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_1_LC_9_7_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance5.Quad_1_LC_9_7_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \QuadInstance5.Quad_1_LC_9_7_7  (
            .in0(N__31248),
            .in1(N__18300),
            .in2(_gnd_net_),
            .in3(N__25735),
            .lcout(dataRead5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38629),
            .ce(),
            .sr(N__35698));
    defparam \QuadInstance7.un1_Quad_cry_0_c_LC_9_8_0 .C_ON=1'b1;
    defparam \QuadInstance7.un1_Quad_cry_0_c_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.un1_Quad_cry_0_c_LC_9_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \QuadInstance7.un1_Quad_cry_0_c_LC_9_8_0  (
            .in0(_gnd_net_),
            .in1(N__21791),
            .in2(N__30776),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(\QuadInstance7.un1_Quad_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNO_0_1_LC_9_8_1 .C_ON=1'b1;
    defparam \QuadInstance7.Quad_RNO_0_1_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNO_0_1_LC_9_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance7.Quad_RNO_0_1_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(N__25842),
            .in2(N__17673),
            .in3(N__17664),
            .lcout(\QuadInstance7.Quad_RNO_0_6_1 ),
            .ltout(),
            .carryin(\QuadInstance7.un1_Quad_cry_0 ),
            .carryout(\QuadInstance7.un1_Quad_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNO_0_2_LC_9_8_2 .C_ON=1'b1;
    defparam \QuadInstance7.Quad_RNO_0_2_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNO_0_2_LC_9_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance7.Quad_RNO_0_2_LC_9_8_2  (
            .in0(_gnd_net_),
            .in1(N__30379),
            .in2(N__17661),
            .in3(N__17652),
            .lcout(\QuadInstance7.Quad_RNO_0_7_2 ),
            .ltout(),
            .carryin(\QuadInstance7.un1_Quad_cry_1 ),
            .carryout(\QuadInstance7.un1_Quad_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNO_0_3_LC_9_8_3 .C_ON=1'b1;
    defparam \QuadInstance7.Quad_RNO_0_3_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNO_0_3_LC_9_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance7.Quad_RNO_0_3_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(N__27841),
            .in2(N__17649),
            .in3(N__17640),
            .lcout(\QuadInstance7.Quad_RNO_0_7_3 ),
            .ltout(),
            .carryin(\QuadInstance7.un1_Quad_cry_2 ),
            .carryout(\QuadInstance7.un1_Quad_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNO_0_4_LC_9_8_4 .C_ON=1'b1;
    defparam \QuadInstance7.Quad_RNO_0_4_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNO_0_4_LC_9_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance7.Quad_RNO_0_4_LC_9_8_4  (
            .in0(_gnd_net_),
            .in1(N__21464),
            .in2(N__17637),
            .in3(N__17628),
            .lcout(\QuadInstance7.Quad_RNO_0_7_4 ),
            .ltout(),
            .carryin(\QuadInstance7.un1_Quad_cry_3 ),
            .carryout(\QuadInstance7.un1_Quad_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNO_0_5_LC_9_8_5 .C_ON=1'b1;
    defparam \QuadInstance7.Quad_RNO_0_5_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNO_0_5_LC_9_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance7.Quad_RNO_0_5_LC_9_8_5  (
            .in0(_gnd_net_),
            .in1(N__36739),
            .in2(N__17625),
            .in3(N__17616),
            .lcout(\QuadInstance7.Quad_RNO_0_7_5 ),
            .ltout(),
            .carryin(\QuadInstance7.un1_Quad_cry_4 ),
            .carryout(\QuadInstance7.un1_Quad_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNO_0_6_LC_9_8_6 .C_ON=1'b1;
    defparam \QuadInstance7.Quad_RNO_0_6_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNO_0_6_LC_9_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance7.Quad_RNO_0_6_LC_9_8_6  (
            .in0(_gnd_net_),
            .in1(N__27700),
            .in2(N__17613),
            .in3(N__17604),
            .lcout(\QuadInstance7.Quad_RNO_0_7_6 ),
            .ltout(),
            .carryin(\QuadInstance7.un1_Quad_cry_5 ),
            .carryout(\QuadInstance7.un1_Quad_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNO_0_7_LC_9_8_7 .C_ON=1'b1;
    defparam \QuadInstance7.Quad_RNO_0_7_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNO_0_7_LC_9_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance7.Quad_RNO_0_7_LC_9_8_7  (
            .in0(_gnd_net_),
            .in1(N__26257),
            .in2(N__17784),
            .in3(N__17775),
            .lcout(\QuadInstance7.Quad_RNO_0_7_7 ),
            .ltout(),
            .carryin(\QuadInstance7.un1_Quad_cry_6 ),
            .carryout(\QuadInstance7.un1_Quad_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNO_0_8_LC_9_9_0 .C_ON=1'b1;
    defparam \QuadInstance7.Quad_RNO_0_8_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNO_0_8_LC_9_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance7.Quad_RNO_0_8_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(N__37612),
            .in2(N__17772),
            .in3(N__17763),
            .lcout(\QuadInstance7.Quad_RNO_0_7_8 ),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(\QuadInstance7.un1_Quad_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNO_0_9_LC_9_9_1 .C_ON=1'b1;
    defparam \QuadInstance7.Quad_RNO_0_9_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNO_0_9_LC_9_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance7.Quad_RNO_0_9_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(N__25387),
            .in2(N__17760),
            .in3(N__17751),
            .lcout(\QuadInstance7.Quad_RNO_0_7_9 ),
            .ltout(),
            .carryin(\QuadInstance7.un1_Quad_cry_8 ),
            .carryout(\QuadInstance7.un1_Quad_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNO_0_10_LC_9_9_2 .C_ON=1'b1;
    defparam \QuadInstance7.Quad_RNO_0_10_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNO_0_10_LC_9_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance7.Quad_RNO_0_10_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(N__34645),
            .in2(N__17748),
            .in3(N__17739),
            .lcout(\QuadInstance7.Quad_RNO_0_7_10 ),
            .ltout(),
            .carryin(\QuadInstance7.un1_Quad_cry_9 ),
            .carryout(\QuadInstance7.un1_Quad_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNO_0_11_LC_9_9_3 .C_ON=1'b1;
    defparam \QuadInstance7.Quad_RNO_0_11_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNO_0_11_LC_9_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance7.Quad_RNO_0_11_LC_9_9_3  (
            .in0(_gnd_net_),
            .in1(N__20875),
            .in2(N__17736),
            .in3(N__17718),
            .lcout(\QuadInstance7.Quad_RNO_0_7_11 ),
            .ltout(),
            .carryin(\QuadInstance7.un1_Quad_cry_10 ),
            .carryout(\QuadInstance7.un1_Quad_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNO_0_12_LC_9_9_4 .C_ON=1'b1;
    defparam \QuadInstance7.Quad_RNO_0_12_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNO_0_12_LC_9_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance7.Quad_RNO_0_12_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(N__22252),
            .in2(N__17715),
            .in3(N__17697),
            .lcout(\QuadInstance7.Quad_RNO_0_7_12 ),
            .ltout(),
            .carryin(\QuadInstance7.un1_Quad_cry_11 ),
            .carryout(\QuadInstance7.un1_Quad_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNO_0_13_LC_9_9_5 .C_ON=1'b1;
    defparam \QuadInstance7.Quad_RNO_0_13_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNO_0_13_LC_9_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance7.Quad_RNO_0_13_LC_9_9_5  (
            .in0(_gnd_net_),
            .in1(N__26108),
            .in2(N__17694),
            .in3(N__17685),
            .lcout(\QuadInstance7.Quad_RNO_0_7_13 ),
            .ltout(),
            .carryin(\QuadInstance7.un1_Quad_cry_12 ),
            .carryout(\QuadInstance7.un1_Quad_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_RNO_0_14_LC_9_9_6 .C_ON=1'b1;
    defparam \QuadInstance7.Quad_RNO_0_14_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \QuadInstance7.Quad_RNO_0_14_LC_9_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance7.Quad_RNO_0_14_LC_9_9_6  (
            .in0(_gnd_net_),
            .in1(N__17682),
            .in2(N__20282),
            .in3(N__17676),
            .lcout(\QuadInstance7.Quad_RNO_0_7_14 ),
            .ltout(),
            .carryin(\QuadInstance7.un1_Quad_cry_13 ),
            .carryout(\QuadInstance7.un1_Quad_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance7.Quad_15_LC_9_9_7 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_15_LC_9_9_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance7.Quad_15_LC_9_9_7 .LUT_INIT=16'b1101000111100010;
    LogicCell40 \QuadInstance7.Quad_15_LC_9_9_7  (
            .in0(N__17835),
            .in1(N__25969),
            .in2(N__31909),
            .in3(N__17826),
            .lcout(dataRead7_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38608),
            .ce(),
            .sr(N__35709));
    defparam \QuadInstance3.Quad_RNIQ30J1_12_LC_9_10_0 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_RNIQ30J1_12_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNIQ30J1_12_LC_9_10_0 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \QuadInstance3.Quad_RNIQ30J1_12_LC_9_10_0  (
            .in0(N__21928),
            .in1(N__19035),
            .in2(N__22332),
            .in3(N__18947),
            .lcout(\QuadInstance3.Quad_RNIQ30J1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_RNIAQAL1_3_LC_9_10_1 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_RNIAQAL1_3_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNIAQAL1_3_LC_9_10_1 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance3.Quad_RNIAQAL1_3_LC_9_10_1  (
            .in0(N__24375),
            .in1(N__21922),
            .in2(N__18971),
            .in3(N__19024),
            .lcout(\QuadInstance3.Quad_RNIAQAL1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_RNIDTAL1_6_LC_9_10_2 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_RNIDTAL1_6_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNIDTAL1_6_LC_9_10_2 .LUT_INIT=16'b1111010100000000;
    LogicCell40 \QuadInstance3.Quad_RNIDTAL1_6_LC_9_10_2  (
            .in0(N__19025),
            .in1(N__28265),
            .in2(N__21969),
            .in3(N__18945),
            .lcout(\QuadInstance3.Quad_RNIDTAL1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_RNICSAL1_5_LC_9_10_3 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_RNICSAL1_5_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNICSAL1_5_LC_9_10_3 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance3.Quad_RNICSAL1_5_LC_9_10_3  (
            .in0(N__23745),
            .in1(N__21923),
            .in2(N__18972),
            .in3(N__19026),
            .lcout(\QuadInstance3.Quad_RNICSAL1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_RNIR40J1_13_LC_9_10_4 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_RNIR40J1_13_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNIR40J1_13_LC_9_10_4 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \QuadInstance3.Quad_RNIR40J1_13_LC_9_10_4  (
            .in0(N__21929),
            .in1(N__19039),
            .in2(N__19938),
            .in3(N__18948),
            .lcout(\QuadInstance3.Quad_RNIR40J1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_RNIP20J1_11_LC_9_10_5 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_RNIP20J1_11_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNIP20J1_11_LC_9_10_5 .LUT_INIT=16'b1000101010001010;
    LogicCell40 \QuadInstance3.Quad_RNIP20J1_11_LC_9_10_5  (
            .in0(N__18946),
            .in1(N__21927),
            .in2(N__19041),
            .in3(N__22422),
            .lcout(\QuadInstance3.Quad_RNIP20J1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwmWrite_fast_1_LC_9_10_6.C_ON=1'b0;
    defparam pwmWrite_fast_1_LC_9_10_6.SEQ_MODE=4'b1000;
    defparam pwmWrite_fast_1_LC_9_10_6.LUT_INIT=16'b0000000000000010;
    LogicCell40 pwmWrite_fast_1_LC_9_10_6 (
            .in0(N__23450),
            .in1(N__33367),
            .in2(N__33671),
            .in3(N__33829),
            .lcout(pwmWrite_fastZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38596),
            .ce(),
            .sr(_gnd_net_));
    defparam pwmWrite_7_LC_9_10_7.C_ON=1'b0;
    defparam pwmWrite_7_LC_9_10_7.SEQ_MODE=4'b1000;
    defparam pwmWrite_7_LC_9_10_7.LUT_INIT=16'b0000100000000000;
    LogicCell40 pwmWrite_7_LC_9_10_7 (
            .in0(N__33828),
            .in1(N__33662),
            .in2(N__33432),
            .in3(N__23449),
            .lcout(pwmWriteZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38596),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.periodCounter_RNIUTF81_13_LC_9_11_0 .C_ON=1'b0;
    defparam \PWMInstance5.periodCounter_RNIUTF81_13_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance5.periodCounter_RNIUTF81_13_LC_9_11_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \PWMInstance5.periodCounter_RNIUTF81_13_LC_9_11_0  (
            .in0(N__17855),
            .in1(N__18173),
            .in2(N__17967),
            .in3(N__17943),
            .lcout(\PWMInstance5.un1_periodCounter12_1_0_a2_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_9_11_1 .C_ON=1'b0;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_9_11_1 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance5.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_9_11_1  (
            .in0(N__17889),
            .in1(N__17854),
            .in2(N__19503),
            .in3(N__17895),
            .lcout(\PWMInstance5.un1_PWMPulseWidthCount_0_I_1_c_RNO_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.PWMPulseWidthCount_esr_0_LC_9_11_2 .C_ON=1'b0;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_0_LC_9_11_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_0_LC_9_11_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \PWMInstance5.PWMPulseWidthCount_esr_0_LC_9_11_2  (
            .in0(N__31374),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PWMInstance5.PWMPulseWidthCountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38588),
            .ce(N__19639),
            .sr(N__35729));
    defparam \PWMInstance5.PWMPulseWidthCount_esr_1_LC_9_11_3 .C_ON=1'b0;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_1_LC_9_11_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_1_LC_9_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance5.PWMPulseWidthCount_esr_1_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31239),
            .lcout(\PWMInstance5.PWMPulseWidthCountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38588),
            .ce(N__19639),
            .sr(N__35729));
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_9_11_4 .C_ON=1'b0;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_9_11_4 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \PWMInstance5.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_9_11_4  (
            .in0(N__17962),
            .in1(N__17871),
            .in2(N__17865),
            .in3(N__19297),
            .lcout(\PWMInstance5.un1_PWMPulseWidthCount_0_I_27_c_RNO_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.PWMPulseWidthCount_esr_6_LC_9_11_5 .C_ON=1'b0;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_6_LC_9_11_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_6_LC_9_11_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \PWMInstance5.PWMPulseWidthCount_esr_6_LC_9_11_5  (
            .in0(N__31087),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PWMInstance5.PWMPulseWidthCountZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38588),
            .ce(N__19639),
            .sr(N__35729));
    defparam \PWMInstance5.PWMPulseWidthCount_esr_7_LC_9_11_6 .C_ON=1'b0;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_7_LC_9_11_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_7_LC_9_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance5.PWMPulseWidthCount_esr_7_LC_9_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29425),
            .lcout(\PWMInstance5.PWMPulseWidthCountZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38588),
            .ce(N__19639),
            .sr(N__35729));
    defparam \PWMInstance5.periodCounter_0_LC_9_12_0 .C_ON=1'b1;
    defparam \PWMInstance5.periodCounter_0_LC_9_12_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.periodCounter_0_LC_9_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance5.periodCounter_0_LC_9_12_0  (
            .in0(_gnd_net_),
            .in1(N__17856),
            .in2(N__19539),
            .in3(N__19538),
            .lcout(\PWMInstance5.periodCounterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_9_12_0_),
            .carryout(\PWMInstance5.un1_periodCounter_2_cry_0 ),
            .clk(N__38577),
            .ce(),
            .sr(N__35307));
    defparam \PWMInstance5.periodCounter_1_LC_9_12_1 .C_ON=1'b1;
    defparam \PWMInstance5.periodCounter_1_LC_9_12_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.periodCounter_1_LC_9_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance5.periodCounter_1_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(N__19502),
            .in2(_gnd_net_),
            .in3(N__17841),
            .lcout(\PWMInstance5.periodCounterZ0Z_1 ),
            .ltout(),
            .carryin(\PWMInstance5.un1_periodCounter_2_cry_0 ),
            .carryout(\PWMInstance5.un1_periodCounter_2_cry_1 ),
            .clk(N__38577),
            .ce(),
            .sr(N__35307));
    defparam \PWMInstance5.periodCounter_2_LC_9_12_2 .C_ON=1'b1;
    defparam \PWMInstance5.periodCounter_2_LC_9_12_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.periodCounter_2_LC_9_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance5.periodCounter_2_LC_9_12_2  (
            .in0(_gnd_net_),
            .in1(N__19257),
            .in2(_gnd_net_),
            .in3(N__17838),
            .lcout(\PWMInstance5.periodCounterZ0Z_2 ),
            .ltout(),
            .carryin(\PWMInstance5.un1_periodCounter_2_cry_1 ),
            .carryout(\PWMInstance5.un1_periodCounter_2_cry_2 ),
            .clk(N__38577),
            .ce(),
            .sr(N__35307));
    defparam \PWMInstance5.periodCounter_3_LC_9_12_3 .C_ON=1'b1;
    defparam \PWMInstance5.periodCounter_3_LC_9_12_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.periodCounter_3_LC_9_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance5.periodCounter_3_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(N__19345),
            .in2(_gnd_net_),
            .in3(N__17976),
            .lcout(\PWMInstance5.periodCounterZ0Z_3 ),
            .ltout(),
            .carryin(\PWMInstance5.un1_periodCounter_2_cry_2 ),
            .carryout(\PWMInstance5.un1_periodCounter_2_cry_3 ),
            .clk(N__38577),
            .ce(),
            .sr(N__35307));
    defparam \PWMInstance5.periodCounter_4_LC_9_12_4 .C_ON=1'b1;
    defparam \PWMInstance5.periodCounter_4_LC_9_12_4 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.periodCounter_4_LC_9_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance5.periodCounter_4_LC_9_12_4  (
            .in0(_gnd_net_),
            .in1(N__19200),
            .in2(_gnd_net_),
            .in3(N__17973),
            .lcout(\PWMInstance5.periodCounterZ0Z_4 ),
            .ltout(),
            .carryin(\PWMInstance5.un1_periodCounter_2_cry_3 ),
            .carryout(\PWMInstance5.un1_periodCounter_2_cry_4 ),
            .clk(N__38577),
            .ce(),
            .sr(N__35307));
    defparam \PWMInstance5.periodCounter_5_LC_9_12_5 .C_ON=1'b1;
    defparam \PWMInstance5.periodCounter_5_LC_9_12_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.periodCounter_5_LC_9_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance5.periodCounter_5_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(N__19393),
            .in2(_gnd_net_),
            .in3(N__17970),
            .lcout(\PWMInstance5.periodCounterZ0Z_5 ),
            .ltout(),
            .carryin(\PWMInstance5.un1_periodCounter_2_cry_4 ),
            .carryout(\PWMInstance5.un1_periodCounter_2_cry_5 ),
            .clk(N__38577),
            .ce(),
            .sr(N__35307));
    defparam \PWMInstance5.periodCounter_6_LC_9_12_6 .C_ON=1'b1;
    defparam \PWMInstance5.periodCounter_6_LC_9_12_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.periodCounter_6_LC_9_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance5.periodCounter_6_LC_9_12_6  (
            .in0(_gnd_net_),
            .in1(N__17966),
            .in2(_gnd_net_),
            .in3(N__17949),
            .lcout(\PWMInstance5.periodCounterZ0Z_6 ),
            .ltout(),
            .carryin(\PWMInstance5.un1_periodCounter_2_cry_5 ),
            .carryout(\PWMInstance5.un1_periodCounter_2_cry_6 ),
            .clk(N__38577),
            .ce(),
            .sr(N__35307));
    defparam \PWMInstance5.periodCounter_7_LC_9_12_7 .C_ON=1'b1;
    defparam \PWMInstance5.periodCounter_7_LC_9_12_7 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.periodCounter_7_LC_9_12_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance5.periodCounter_7_LC_9_12_7  (
            .in0(N__19451),
            .in1(N__19298),
            .in2(_gnd_net_),
            .in3(N__17946),
            .lcout(\PWMInstance5.periodCounterZ0Z_7 ),
            .ltout(),
            .carryin(\PWMInstance5.un1_periodCounter_2_cry_6 ),
            .carryout(\PWMInstance5.un1_periodCounter_2_cry_7 ),
            .clk(N__38577),
            .ce(),
            .sr(N__35307));
    defparam \PWMInstance5.periodCounter_8_LC_9_13_0 .C_ON=1'b1;
    defparam \PWMInstance5.periodCounter_8_LC_9_13_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.periodCounter_8_LC_9_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance5.periodCounter_8_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(N__17941),
            .in2(_gnd_net_),
            .in3(N__17919),
            .lcout(\PWMInstance5.periodCounterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_9_13_0_),
            .carryout(\PWMInstance5.un1_periodCounter_2_cry_8 ),
            .clk(N__38567),
            .ce(),
            .sr(N__35306));
    defparam \PWMInstance5.periodCounter_9_LC_9_13_1 .C_ON=1'b1;
    defparam \PWMInstance5.periodCounter_9_LC_9_13_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.periodCounter_9_LC_9_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance5.periodCounter_9_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(N__19415),
            .in2(_gnd_net_),
            .in3(N__17916),
            .lcout(\PWMInstance5.periodCounterZ0Z_9 ),
            .ltout(),
            .carryin(\PWMInstance5.un1_periodCounter_2_cry_8 ),
            .carryout(\PWMInstance5.un1_periodCounter_2_cry_9 ),
            .clk(N__38567),
            .ce(),
            .sr(N__35306));
    defparam \PWMInstance5.periodCounter_10_LC_9_13_2 .C_ON=1'b1;
    defparam \PWMInstance5.periodCounter_10_LC_9_13_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.periodCounter_10_LC_9_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance5.periodCounter_10_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(N__19173),
            .in2(_gnd_net_),
            .in3(N__17913),
            .lcout(\PWMInstance5.periodCounterZ0Z_10 ),
            .ltout(),
            .carryin(\PWMInstance5.un1_periodCounter_2_cry_9 ),
            .carryout(\PWMInstance5.un1_periodCounter_2_cry_10 ),
            .clk(N__38567),
            .ce(),
            .sr(N__35306));
    defparam \PWMInstance5.periodCounter_11_LC_9_13_3 .C_ON=1'b1;
    defparam \PWMInstance5.periodCounter_11_LC_9_13_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.periodCounter_11_LC_9_13_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance5.periodCounter_11_LC_9_13_3  (
            .in0(N__19453),
            .in1(N__19369),
            .in2(_gnd_net_),
            .in3(N__17910),
            .lcout(\PWMInstance5.periodCounterZ0Z_11 ),
            .ltout(),
            .carryin(\PWMInstance5.un1_periodCounter_2_cry_10 ),
            .carryout(\PWMInstance5.un1_periodCounter_2_cry_11 ),
            .clk(N__38567),
            .ce(),
            .sr(N__35306));
    defparam \PWMInstance5.periodCounter_12_LC_9_13_4 .C_ON=1'b1;
    defparam \PWMInstance5.periodCounter_12_LC_9_13_4 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.periodCounter_12_LC_9_13_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance5.periodCounter_12_LC_9_13_4  (
            .in0(N__19450),
            .in1(N__19221),
            .in2(_gnd_net_),
            .in3(N__18180),
            .lcout(\PWMInstance5.periodCounterZ0Z_12 ),
            .ltout(),
            .carryin(\PWMInstance5.un1_periodCounter_2_cry_11 ),
            .carryout(\PWMInstance5.un1_periodCounter_2_cry_12 ),
            .clk(N__38567),
            .ce(),
            .sr(N__35306));
    defparam \PWMInstance5.periodCounter_13_LC_9_13_5 .C_ON=1'b1;
    defparam \PWMInstance5.periodCounter_13_LC_9_13_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.periodCounter_13_LC_9_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance5.periodCounter_13_LC_9_13_5  (
            .in0(N__19454),
            .in1(N__18172),
            .in2(_gnd_net_),
            .in3(N__18153),
            .lcout(\PWMInstance5.periodCounterZ0Z_13 ),
            .ltout(),
            .carryin(\PWMInstance5.un1_periodCounter_2_cry_12 ),
            .carryout(\PWMInstance5.un1_periodCounter_2_cry_13 ),
            .clk(N__38567),
            .ce(),
            .sr(N__35306));
    defparam \PWMInstance5.periodCounter_14_LC_9_13_6 .C_ON=1'b1;
    defparam \PWMInstance5.periodCounter_14_LC_9_13_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.periodCounter_14_LC_9_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance5.periodCounter_14_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(N__19239),
            .in2(_gnd_net_),
            .in3(N__18150),
            .lcout(\PWMInstance5.periodCounterZ0Z_14 ),
            .ltout(),
            .carryin(\PWMInstance5.un1_periodCounter_2_cry_13 ),
            .carryout(\PWMInstance5.un1_periodCounter_2_cry_14 ),
            .clk(N__38567),
            .ce(),
            .sr(N__35306));
    defparam \PWMInstance5.periodCounter_15_LC_9_13_7 .C_ON=1'b1;
    defparam \PWMInstance5.periodCounter_15_LC_9_13_7 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.periodCounter_15_LC_9_13_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance5.periodCounter_15_LC_9_13_7  (
            .in0(_gnd_net_),
            .in1(N__19523),
            .in2(_gnd_net_),
            .in3(N__18147),
            .lcout(\PWMInstance5.periodCounterZ0Z_15 ),
            .ltout(),
            .carryin(\PWMInstance5.un1_periodCounter_2_cry_14 ),
            .carryout(\PWMInstance5.un1_periodCounter_2_cry_15 ),
            .clk(N__38567),
            .ce(),
            .sr(N__35306));
    defparam \PWMInstance5.periodCounter_16_LC_9_14_0 .C_ON=1'b0;
    defparam \PWMInstance5.periodCounter_16_LC_9_14_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.periodCounter_16_LC_9_14_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance5.periodCounter_16_LC_9_14_0  (
            .in0(N__19452),
            .in1(N__19317),
            .in2(_gnd_net_),
            .in3(N__18144),
            .lcout(\PWMInstance5.periodCounterZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38561),
            .ce(),
            .sr(N__35304));
    defparam \PWMInstance0.periodCounter_RNIA4GO1_13_LC_9_15_0 .C_ON=1'b0;
    defparam \PWMInstance0.periodCounter_RNIA4GO1_13_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance0.periodCounter_RNIA4GO1_13_LC_9_15_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \PWMInstance0.periodCounter_RNIA4GO1_13_LC_9_15_0  (
            .in0(N__18141),
            .in1(N__18110),
            .in2(N__18078),
            .in3(N__18036),
            .lcout(\PWMInstance0.un1_periodCounter12_1_0_a2_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_9_15_1 .C_ON=1'b0;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance0.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_9_15_1 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \PWMInstance0.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_9_15_1  (
            .in0(N__18035),
            .in1(N__18267),
            .in2(N__18015),
            .in3(N__17982),
            .lcout(\PWMInstance0.un1_PWMPulseWidthCount_0_I_1_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance0.PWMPulseWidthCount_esr_0_LC_9_15_2 .C_ON=1'b0;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_0_LC_9_15_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_0_LC_9_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance0.PWMPulseWidthCount_esr_0_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31422),
            .lcout(\PWMInstance0.PWMPulseWidthCountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38554),
            .ce(N__18248),
            .sr(N__35756));
    defparam \PWMInstance0.PWMPulseWidthCount_esr_1_LC_9_15_3 .C_ON=1'b0;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_1_LC_9_15_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_1_LC_9_15_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \PWMInstance0.PWMPulseWidthCount_esr_1_LC_9_15_3  (
            .in0(N__31264),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PWMInstance0.PWMPulseWidthCountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38554),
            .ce(N__18248),
            .sr(N__35756));
    defparam \PWMInstance0.PWMPulseWidthCount_esr_7_LC_9_15_6 .C_ON=1'b0;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_7_LC_9_15_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance0.PWMPulseWidthCount_esr_7_LC_9_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance0.PWMPulseWidthCount_esr_7_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29456),
            .lcout(\PWMInstance0.PWMPulseWidthCountZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38554),
            .ce(N__18248),
            .sr(N__35756));
    defparam \PWMInstance5.PWMPulseWidthCount_esr_13_LC_9_16_4 .C_ON=1'b0;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_13_LC_9_16_4 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_13_LC_9_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance5.PWMPulseWidthCount_esr_13_LC_9_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28726),
            .lcout(\PWMInstance5.PWMPulseWidthCountZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38549),
            .ce(N__19649),
            .sr(N__35759));
    defparam \QuadInstance5.delayedCh_B_0_LC_10_1_7 .C_ON=1'b0;
    defparam \QuadInstance5.delayedCh_B_0_LC_10_1_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance5.delayedCh_B_0_LC_10_1_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance5.delayedCh_B_0_LC_10_1_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18201),
            .lcout(\QuadInstance5.delayedCh_BZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38688),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.delayedCh_A_2_LC_10_4_1 .C_ON=1'b0;
    defparam \QuadInstance5.delayedCh_A_2_LC_10_4_1 .SEQ_MODE=4'b1000;
    defparam \QuadInstance5.delayedCh_A_2_LC_10_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance5.delayedCh_A_2_LC_10_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18435),
            .lcout(\QuadInstance5.delayedCh_AZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38661),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.delayedCh_B_1_LC_10_4_5 .C_ON=1'b0;
    defparam \QuadInstance5.delayedCh_B_1_LC_10_4_5 .SEQ_MODE=4'b1000;
    defparam \QuadInstance5.delayedCh_B_1_LC_10_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance5.delayedCh_B_1_LC_10_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18189),
            .lcout(\QuadInstance5.delayedCh_BZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38661),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.delayedCh_B_2_LC_10_4_6 .C_ON=1'b0;
    defparam \QuadInstance5.delayedCh_B_2_LC_10_4_6 .SEQ_MODE=4'b1000;
    defparam \QuadInstance5.delayedCh_B_2_LC_10_4_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance5.delayedCh_B_2_LC_10_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18447),
            .lcout(\QuadInstance5.delayedCh_BZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38661),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_RNO_0_15_LC_10_5_0 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_RNO_0_15_LC_10_5_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNO_0_15_LC_10_5_0 .LUT_INIT=16'b0100101111110000;
    LogicCell40 \QuadInstance4.Quad_RNO_0_15_LC_10_5_0  (
            .in0(N__29663),
            .in1(N__27354),
            .in2(N__25224),
            .in3(N__27452),
            .lcout(\QuadInstance4.un1_Quad_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_0_LC_10_5_1 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_0_LC_10_5_1 .SEQ_MODE=4'b1000;
    defparam \QuadInstance4.Quad_0_LC_10_5_1 .LUT_INIT=16'b1111000001100110;
    LogicCell40 \QuadInstance4.Quad_0_LC_10_5_1  (
            .in0(N__27453),
            .in1(N__30268),
            .in2(N__31440),
            .in3(N__29664),
            .lcout(dataRead4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38649),
            .ce(),
            .sr(N__35689));
    defparam \QuadInstance0.Quad_0_LC_10_5_2 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_0_LC_10_5_2 .SEQ_MODE=4'b1000;
    defparam \QuadInstance0.Quad_0_LC_10_5_2 .LUT_INIT=16'b1101000111100010;
    LogicCell40 \QuadInstance0.Quad_0_LC_10_5_2  (
            .in0(N__30299),
            .in1(N__33127),
            .in2(N__31438),
            .in3(N__34089),
            .lcout(dataRead0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38649),
            .ce(),
            .sr(N__35689));
    defparam \QuadInstance2.Quad_0_LC_10_5_3 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_0_LC_10_5_3 .SEQ_MODE=4'b1000;
    defparam \QuadInstance2.Quad_0_LC_10_5_3 .LUT_INIT=16'b1111011000000110;
    LogicCell40 \QuadInstance2.Quad_0_LC_10_5_3  (
            .in0(N__18534),
            .in1(N__30838),
            .in2(N__22190),
            .in3(N__31429),
            .lcout(dataRead2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38649),
            .ce(),
            .sr(N__35689));
    defparam \QuadInstance5.delayedCh_A_RNI0UF71_2_LC_10_5_4 .C_ON=1'b0;
    defparam \QuadInstance5.delayedCh_A_RNI0UF71_2_LC_10_5_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.delayedCh_A_RNI0UF71_2_LC_10_5_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \QuadInstance5.delayedCh_A_RNI0UF71_2_LC_10_5_4  (
            .in0(N__18446),
            .in1(N__18434),
            .in2(N__18417),
            .in3(N__18408),
            .lcout(\QuadInstance5.count_enable ),
            .ltout(\QuadInstance5.count_enable_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_0_LC_10_5_5 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_0_LC_10_5_5 .SEQ_MODE=4'b1000;
    defparam \QuadInstance5.Quad_0_LC_10_5_5 .LUT_INIT=16'b1011111000010100;
    LogicCell40 \QuadInstance5.Quad_0_LC_10_5_5  (
            .in0(N__25778),
            .in1(N__30907),
            .in2(N__18396),
            .in3(N__31430),
            .lcout(dataRead5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38649),
            .ce(),
            .sr(N__35689));
    defparam \QuadInstance3.Quad_0_LC_10_5_6 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_0_LC_10_5_6 .SEQ_MODE=4'b1000;
    defparam \QuadInstance3.Quad_0_LC_10_5_6 .LUT_INIT=16'b1011000111100100;
    LogicCell40 \QuadInstance3.Quad_0_LC_10_5_6  (
            .in0(N__22008),
            .in1(N__30877),
            .in2(N__31439),
            .in3(N__18978),
            .lcout(dataRead3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38649),
            .ce(),
            .sr(N__35689));
    defparam \QuadInstance5.un1_Quad_cry_0_c_LC_10_6_0 .C_ON=1'b1;
    defparam \QuadInstance5.un1_Quad_cry_0_c_LC_10_6_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.un1_Quad_cry_0_c_LC_10_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \QuadInstance5.un1_Quad_cry_0_c_LC_10_6_0  (
            .in0(_gnd_net_),
            .in1(N__18369),
            .in2(N__30908),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_6_0_),
            .carryout(\QuadInstance5.un1_Quad_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNO_0_1_LC_10_6_1 .C_ON=1'b1;
    defparam \QuadInstance5.Quad_RNO_0_1_LC_10_6_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNO_0_1_LC_10_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance5.Quad_RNO_0_1_LC_10_6_1  (
            .in0(_gnd_net_),
            .in1(N__23854),
            .in2(N__18309),
            .in3(N__18294),
            .lcout(\QuadInstance5.Quad_RNO_0_4_1 ),
            .ltout(),
            .carryin(\QuadInstance5.un1_Quad_cry_0 ),
            .carryout(\QuadInstance5.un1_Quad_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNO_0_2_LC_10_6_2 .C_ON=1'b1;
    defparam \QuadInstance5.Quad_RNO_0_2_LC_10_6_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNO_0_2_LC_10_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance5.Quad_RNO_0_2_LC_10_6_2  (
            .in0(_gnd_net_),
            .in1(N__30526),
            .in2(N__18291),
            .in3(N__18282),
            .lcout(\QuadInstance5.Quad_RNO_0_5_2 ),
            .ltout(),
            .carryin(\QuadInstance5.un1_Quad_cry_1 ),
            .carryout(\QuadInstance5.un1_Quad_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNO_0_3_LC_10_6_3 .C_ON=1'b1;
    defparam \QuadInstance5.Quad_RNO_0_3_LC_10_6_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNO_0_3_LC_10_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance5.Quad_RNO_0_3_LC_10_6_3  (
            .in0(_gnd_net_),
            .in1(N__27917),
            .in2(N__18279),
            .in3(N__18270),
            .lcout(\QuadInstance5.Quad_RNO_0_5_3 ),
            .ltout(),
            .carryin(\QuadInstance5.un1_Quad_cry_2 ),
            .carryout(\QuadInstance5.un1_Quad_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNO_0_4_LC_10_6_4 .C_ON=1'b1;
    defparam \QuadInstance5.Quad_RNO_0_4_LC_10_6_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNO_0_4_LC_10_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance5.Quad_RNO_0_4_LC_10_6_4  (
            .in0(_gnd_net_),
            .in1(N__21316),
            .in2(N__18648),
            .in3(N__18639),
            .lcout(\QuadInstance5.Quad_RNO_0_5_4 ),
            .ltout(),
            .carryin(\QuadInstance5.un1_Quad_cry_3 ),
            .carryout(\QuadInstance5.un1_Quad_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNO_0_5_LC_10_6_5 .C_ON=1'b1;
    defparam \QuadInstance5.Quad_RNO_0_5_LC_10_6_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNO_0_5_LC_10_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance5.Quad_RNO_0_5_LC_10_6_5  (
            .in0(_gnd_net_),
            .in1(N__36872),
            .in2(N__18636),
            .in3(N__18627),
            .lcout(\QuadInstance5.Quad_RNO_0_5_5 ),
            .ltout(),
            .carryin(\QuadInstance5.un1_Quad_cry_4 ),
            .carryout(\QuadInstance5.un1_Quad_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNO_0_6_LC_10_6_6 .C_ON=1'b1;
    defparam \QuadInstance5.Quad_RNO_0_6_LC_10_6_6 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNO_0_6_LC_10_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance5.Quad_RNO_0_6_LC_10_6_6  (
            .in0(_gnd_net_),
            .in1(N__25267),
            .in2(N__18624),
            .in3(N__18615),
            .lcout(\QuadInstance5.Quad_RNO_0_5_6 ),
            .ltout(),
            .carryin(\QuadInstance5.un1_Quad_cry_5 ),
            .carryout(\QuadInstance5.un1_Quad_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNO_0_7_LC_10_6_7 .C_ON=1'b1;
    defparam \QuadInstance5.Quad_RNO_0_7_LC_10_6_7 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNO_0_7_LC_10_6_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance5.Quad_RNO_0_7_LC_10_6_7  (
            .in0(_gnd_net_),
            .in1(N__18612),
            .in2(N__25597),
            .in3(N__18606),
            .lcout(\QuadInstance5.Quad_RNO_0_5_7 ),
            .ltout(),
            .carryin(\QuadInstance5.un1_Quad_cry_6 ),
            .carryout(\QuadInstance5.un1_Quad_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNO_0_8_LC_10_7_0 .C_ON=1'b1;
    defparam \QuadInstance5.Quad_RNO_0_8_LC_10_7_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNO_0_8_LC_10_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance5.Quad_RNO_0_8_LC_10_7_0  (
            .in0(_gnd_net_),
            .in1(N__36973),
            .in2(N__18603),
            .in3(N__18594),
            .lcout(\QuadInstance5.Quad_RNO_0_5_8 ),
            .ltout(),
            .carryin(bfn_10_7_0_),
            .carryout(\QuadInstance5.un1_Quad_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNO_0_9_LC_10_7_1 .C_ON=1'b1;
    defparam \QuadInstance5.Quad_RNO_0_9_LC_10_7_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNO_0_9_LC_10_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance5.Quad_RNO_0_9_LC_10_7_1  (
            .in0(_gnd_net_),
            .in1(N__25507),
            .in2(N__18591),
            .in3(N__18579),
            .lcout(\QuadInstance5.Quad_RNO_0_5_9 ),
            .ltout(),
            .carryin(\QuadInstance5.un1_Quad_cry_8 ),
            .carryout(\QuadInstance5.un1_Quad_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNO_0_10_LC_10_7_2 .C_ON=1'b1;
    defparam \QuadInstance5.Quad_RNO_0_10_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNO_0_10_LC_10_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance5.Quad_RNO_0_10_LC_10_7_2  (
            .in0(_gnd_net_),
            .in1(N__35008),
            .in2(N__18576),
            .in3(N__18567),
            .lcout(\QuadInstance5.Quad_RNO_0_5_10 ),
            .ltout(),
            .carryin(\QuadInstance5.un1_Quad_cry_9 ),
            .carryout(\QuadInstance5.un1_Quad_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNO_0_11_LC_10_7_3 .C_ON=1'b1;
    defparam \QuadInstance5.Quad_RNO_0_11_LC_10_7_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNO_0_11_LC_10_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance5.Quad_RNO_0_11_LC_10_7_3  (
            .in0(_gnd_net_),
            .in1(N__20101),
            .in2(N__18564),
            .in3(N__18555),
            .lcout(\QuadInstance5.Quad_RNO_0_5_11 ),
            .ltout(),
            .carryin(\QuadInstance5.un1_Quad_cry_10 ),
            .carryout(\QuadInstance5.un1_Quad_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNO_0_12_LC_10_7_4 .C_ON=1'b1;
    defparam \QuadInstance5.Quad_RNO_0_12_LC_10_7_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNO_0_12_LC_10_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance5.Quad_RNO_0_12_LC_10_7_4  (
            .in0(_gnd_net_),
            .in1(N__22378),
            .in2(N__18552),
            .in3(N__18537),
            .lcout(\QuadInstance5.Quad_RNO_0_5_12 ),
            .ltout(),
            .carryin(\QuadInstance5.un1_Quad_cry_11 ),
            .carryout(\QuadInstance5.un1_Quad_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNO_0_13_LC_10_7_5 .C_ON=1'b1;
    defparam \QuadInstance5.Quad_RNO_0_13_LC_10_7_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNO_0_13_LC_10_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance5.Quad_RNO_0_13_LC_10_7_5  (
            .in0(_gnd_net_),
            .in1(N__18711),
            .in2(N__20012),
            .in3(N__18699),
            .lcout(\QuadInstance5.Quad_RNO_0_5_13 ),
            .ltout(),
            .carryin(\QuadInstance5.un1_Quad_cry_12 ),
            .carryout(\QuadInstance5.un1_Quad_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_RNO_0_14_LC_10_7_6 .C_ON=1'b1;
    defparam \QuadInstance5.Quad_RNO_0_14_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \QuadInstance5.Quad_RNO_0_14_LC_10_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance5.Quad_RNO_0_14_LC_10_7_6  (
            .in0(_gnd_net_),
            .in1(N__18696),
            .in2(N__28226),
            .in3(N__18684),
            .lcout(\QuadInstance5.Quad_RNO_0_5_14 ),
            .ltout(),
            .carryin(\QuadInstance5.un1_Quad_cry_13 ),
            .carryout(\QuadInstance5.un1_Quad_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance5.Quad_15_LC_10_7_7 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_15_LC_10_7_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance5.Quad_15_LC_10_7_7 .LUT_INIT=16'b1101000111100010;
    LogicCell40 \QuadInstance5.Quad_15_LC_10_7_7  (
            .in0(N__18681),
            .in1(N__25756),
            .in2(N__31919),
            .in3(N__18675),
            .lcout(dataRead5_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38630),
            .ce(),
            .sr(N__35699));
    defparam \QuadInstance3.un1_Quad_cry_0_c_LC_10_8_0 .C_ON=1'b1;
    defparam \QuadInstance3.un1_Quad_cry_0_c_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.un1_Quad_cry_0_c_LC_10_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \QuadInstance3.un1_Quad_cry_0_c_LC_10_8_0  (
            .in0(_gnd_net_),
            .in1(N__18976),
            .in2(N__30878),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_8_0_),
            .carryout(\QuadInstance3.un1_Quad_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_RNO_0_1_LC_10_8_1 .C_ON=1'b1;
    defparam \QuadInstance3.Quad_RNO_0_1_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNO_0_1_LC_10_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance3.Quad_RNO_0_1_LC_10_8_1  (
            .in0(_gnd_net_),
            .in1(N__23807),
            .in2(N__18843),
            .in3(N__18672),
            .lcout(\QuadInstance3.Quad_RNO_0_2_1 ),
            .ltout(),
            .carryin(\QuadInstance3.un1_Quad_cry_0 ),
            .carryout(\QuadInstance3.un1_Quad_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_RNO_0_2_LC_10_8_2 .C_ON=1'b1;
    defparam \QuadInstance3.Quad_RNO_0_2_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNO_0_2_LC_10_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance3.Quad_RNO_0_2_LC_10_8_2  (
            .in0(_gnd_net_),
            .in1(N__30418),
            .in2(N__18828),
            .in3(N__18669),
            .lcout(\QuadInstance3.Quad_RNO_0_3_2 ),
            .ltout(),
            .carryin(\QuadInstance3.un1_Quad_cry_1 ),
            .carryout(\QuadInstance3.un1_Quad_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_RNO_0_3_LC_10_8_3 .C_ON=1'b1;
    defparam \QuadInstance3.Quad_RNO_0_3_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNO_0_3_LC_10_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance3.Quad_RNO_0_3_LC_10_8_3  (
            .in0(_gnd_net_),
            .in1(N__24367),
            .in2(N__18666),
            .in3(N__18654),
            .lcout(\QuadInstance3.Quad_RNO_0_3_3 ),
            .ltout(),
            .carryin(\QuadInstance3.un1_Quad_cry_2 ),
            .carryout(\QuadInstance3.un1_Quad_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_RNO_0_4_LC_10_8_4 .C_ON=1'b1;
    defparam \QuadInstance3.Quad_RNO_0_4_LC_10_8_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNO_0_4_LC_10_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance3.Quad_RNO_0_4_LC_10_8_4  (
            .in0(_gnd_net_),
            .in1(N__19107),
            .in2(N__21845),
            .in3(N__18651),
            .lcout(\QuadInstance3.Quad_RNO_0_3_4 ),
            .ltout(),
            .carryin(\QuadInstance3.un1_Quad_cry_3 ),
            .carryout(\QuadInstance3.un1_Quad_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_RNO_0_5_LC_10_8_5 .C_ON=1'b1;
    defparam \QuadInstance3.Quad_RNO_0_5_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNO_0_5_LC_10_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance3.Quad_RNO_0_5_LC_10_8_5  (
            .in0(_gnd_net_),
            .in1(N__23741),
            .in2(N__18789),
            .in3(N__18777),
            .lcout(\QuadInstance3.Quad_RNO_0_3_5 ),
            .ltout(),
            .carryin(\QuadInstance3.un1_Quad_cry_4 ),
            .carryout(\QuadInstance3.un1_Quad_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_RNO_0_6_LC_10_8_6 .C_ON=1'b1;
    defparam \QuadInstance3.Quad_RNO_0_6_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNO_0_6_LC_10_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance3.Quad_RNO_0_6_LC_10_8_6  (
            .in0(_gnd_net_),
            .in1(N__28258),
            .in2(N__18774),
            .in3(N__18762),
            .lcout(\QuadInstance3.Quad_RNO_0_3_6 ),
            .ltout(),
            .carryin(\QuadInstance3.un1_Quad_cry_5 ),
            .carryout(\QuadInstance3.un1_Quad_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_RNO_0_7_LC_10_8_7 .C_ON=1'b1;
    defparam \QuadInstance3.Quad_RNO_0_7_LC_10_8_7 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNO_0_7_LC_10_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance3.Quad_RNO_0_7_LC_10_8_7  (
            .in0(_gnd_net_),
            .in1(N__26329),
            .in2(N__19053),
            .in3(N__18759),
            .lcout(\QuadInstance3.Quad_RNO_0_3_7 ),
            .ltout(),
            .carryin(\QuadInstance3.un1_Quad_cry_6 ),
            .carryout(\QuadInstance3.un1_Quad_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_RNO_0_8_LC_10_9_0 .C_ON=1'b1;
    defparam \QuadInstance3.Quad_RNO_0_8_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNO_0_8_LC_10_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance3.Quad_RNO_0_8_LC_10_9_0  (
            .in0(_gnd_net_),
            .in1(N__30661),
            .in2(N__18807),
            .in3(N__18756),
            .lcout(\QuadInstance3.Quad_RNO_0_3_8 ),
            .ltout(),
            .carryin(bfn_10_9_0_),
            .carryout(\QuadInstance3.un1_Quad_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_RNO_0_9_LC_10_9_1 .C_ON=1'b1;
    defparam \QuadInstance3.Quad_RNO_0_9_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNO_0_9_LC_10_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance3.Quad_RNO_0_9_LC_10_9_1  (
            .in0(_gnd_net_),
            .in1(N__25480),
            .in2(N__18798),
            .in3(N__18753),
            .lcout(\QuadInstance3.Quad_RNO_0_3_9 ),
            .ltout(),
            .carryin(\QuadInstance3.un1_Quad_cry_8 ),
            .carryout(\QuadInstance3.un1_Quad_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_RNO_0_10_LC_10_9_2 .C_ON=1'b1;
    defparam \QuadInstance3.Quad_RNO_0_10_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNO_0_10_LC_10_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance3.Quad_RNO_0_10_LC_10_9_2  (
            .in0(_gnd_net_),
            .in1(N__34789),
            .in2(N__18816),
            .in3(N__18750),
            .lcout(\QuadInstance3.Quad_RNO_0_3_10 ),
            .ltout(),
            .carryin(\QuadInstance3.un1_Quad_cry_9 ),
            .carryout(\QuadInstance3.un1_Quad_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_RNO_0_11_LC_10_9_3 .C_ON=1'b1;
    defparam \QuadInstance3.Quad_RNO_0_11_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNO_0_11_LC_10_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance3.Quad_RNO_0_11_LC_10_9_3  (
            .in0(_gnd_net_),
            .in1(N__22414),
            .in2(N__18747),
            .in3(N__18738),
            .lcout(\QuadInstance3.Quad_RNO_0_3_11 ),
            .ltout(),
            .carryin(\QuadInstance3.un1_Quad_cry_10 ),
            .carryout(\QuadInstance3.un1_Quad_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_RNO_0_12_LC_10_9_4 .C_ON=1'b1;
    defparam \QuadInstance3.Quad_RNO_0_12_LC_10_9_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNO_0_12_LC_10_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance3.Quad_RNO_0_12_LC_10_9_4  (
            .in0(_gnd_net_),
            .in1(N__22315),
            .in2(N__18735),
            .in3(N__18726),
            .lcout(\QuadInstance3.Quad_RNO_0_3_12 ),
            .ltout(),
            .carryin(\QuadInstance3.un1_Quad_cry_11 ),
            .carryout(\QuadInstance3.un1_Quad_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_RNO_0_13_LC_10_9_5 .C_ON=1'b1;
    defparam \QuadInstance3.Quad_RNO_0_13_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNO_0_13_LC_10_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance3.Quad_RNO_0_13_LC_10_9_5  (
            .in0(_gnd_net_),
            .in1(N__19928),
            .in2(N__18723),
            .in3(N__18714),
            .lcout(\QuadInstance3.Quad_RNO_0_3_13 ),
            .ltout(),
            .carryin(\QuadInstance3.un1_Quad_cry_12 ),
            .carryout(\QuadInstance3.un1_Quad_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_RNO_0_14_LC_10_9_6 .C_ON=1'b1;
    defparam \QuadInstance3.Quad_RNO_0_14_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNO_0_14_LC_10_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance3.Quad_RNO_0_14_LC_10_9_6  (
            .in0(_gnd_net_),
            .in1(N__19098),
            .in2(N__20072),
            .in3(N__18852),
            .lcout(\QuadInstance3.Quad_RNO_0_3_14 ),
            .ltout(),
            .carryin(\QuadInstance3.un1_Quad_cry_13 ),
            .carryout(\QuadInstance3.un1_Quad_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_15_LC_10_9_7 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_15_LC_10_9_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance3.Quad_15_LC_10_9_7 .LUT_INIT=16'b1101000111100010;
    LogicCell40 \QuadInstance3.Quad_15_LC_10_9_7  (
            .in0(N__18888),
            .in1(N__21985),
            .in2(N__31908),
            .in3(N__18849),
            .lcout(dataRead3_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38609),
            .ce(),
            .sr(N__35713));
    defparam \QuadInstance3.delayedCh_A_RNIO54L_2_LC_10_10_0 .C_ON=1'b0;
    defparam \QuadInstance3.delayedCh_A_RNIO54L_2_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.delayedCh_A_RNIO54L_2_LC_10_10_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \QuadInstance3.delayedCh_A_RNIO54L_2_LC_10_10_0  (
            .in0(N__19074),
            .in1(N__19067),
            .in2(N__19089),
            .in3(N__18863),
            .lcout(\QuadInstance3.count_enable ),
            .ltout(\QuadInstance3.count_enable_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_RNI8OAL1_1_LC_10_10_1 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_RNI8OAL1_1_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNI8OAL1_1_LC_10_10_1 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance3.Quad_RNI8OAL1_1_LC_10_10_1  (
            .in0(N__23811),
            .in1(N__21917),
            .in2(N__18846),
            .in3(N__19022),
            .lcout(\QuadInstance3.Quad_RNI8OAL1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.delayedCh_B_RNIQUMH_2_LC_10_10_2 .C_ON=1'b0;
    defparam \QuadInstance3.delayedCh_B_RNIQUMH_2_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.delayedCh_B_RNIQUMH_2_LC_10_10_2 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \QuadInstance3.delayedCh_B_RNIQUMH_2_LC_10_10_2  (
            .in0(N__34501),
            .in1(_gnd_net_),
            .in2(N__19088),
            .in3(N__19066),
            .lcout(\QuadInstance3.un1_count_enable_i_a2_0_1 ),
            .ltout(\QuadInstance3.un1_count_enable_i_a2_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_RNI9PAL1_2_LC_10_10_3 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_RNI9PAL1_2_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNI9PAL1_2_LC_10_10_3 .LUT_INIT=16'b1100111100000000;
    LogicCell40 \QuadInstance3.Quad_RNI9PAL1_2_LC_10_10_3  (
            .in0(N__30422),
            .in1(N__21918),
            .in2(N__18831),
            .in3(N__18949),
            .lcout(\QuadInstance3.Quad_RNI9PAL1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_RNIO10J1_10_LC_10_10_4 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_RNIO10J1_10_LC_10_10_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNIO10J1_10_LC_10_10_4 .LUT_INIT=16'b1011000010110000;
    LogicCell40 \QuadInstance3.Quad_RNIO10J1_10_LC_10_10_4  (
            .in0(N__21921),
            .in1(N__19034),
            .in2(N__18974),
            .in3(N__34803),
            .lcout(\QuadInstance3.Quad_RNIO10J1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_RNIFVAL1_8_LC_10_10_5 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_RNIFVAL1_8_LC_10_10_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNIFVAL1_8_LC_10_10_5 .LUT_INIT=16'b1100111100000000;
    LogicCell40 \QuadInstance3.Quad_RNIFVAL1_8_LC_10_10_5  (
            .in0(N__30668),
            .in1(N__21919),
            .in2(N__19040),
            .in3(N__18954),
            .lcout(\QuadInstance3.Quad_RNIFVAL1Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_RNIG0BL1_9_LC_10_10_6 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_RNIG0BL1_9_LC_10_10_6 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNIG0BL1_9_LC_10_10_6 .LUT_INIT=16'b1011000010110000;
    LogicCell40 \QuadInstance3.Quad_RNIG0BL1_9_LC_10_10_6  (
            .in0(N__21920),
            .in1(N__19030),
            .in2(N__18973),
            .in3(N__25481),
            .lcout(\QuadInstance3.Quad_RNIG0BL1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_RNIBRAL1_4_LC_10_10_7 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_RNIBRAL1_4_LC_10_10_7 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNIBRAL1_4_LC_10_10_7 .LUT_INIT=16'b1100000011001100;
    LogicCell40 \QuadInstance3.Quad_RNIBRAL1_4_LC_10_10_7  (
            .in0(N__21846),
            .in1(N__18950),
            .in2(N__21970),
            .in3(N__19023),
            .lcout(\QuadInstance3.Quad_RNIBRAL1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_RNIS50J1_14_LC_10_11_0 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_RNIS50J1_14_LC_10_11_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNIS50J1_14_LC_10_11_0 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \QuadInstance3.Quad_RNIS50J1_14_LC_10_11_0  (
            .in0(N__21934),
            .in1(N__18964),
            .in2(N__20079),
            .in3(N__19028),
            .lcout(\QuadInstance3.Quad_RNIS50J1Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.delayedCh_B_2_LC_10_11_1 .C_ON=1'b0;
    defparam \QuadInstance3.delayedCh_B_2_LC_10_11_1 .SEQ_MODE=4'b1000;
    defparam \QuadInstance3.delayedCh_B_2_LC_10_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance3.delayedCh_B_2_LC_10_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18864),
            .lcout(\QuadInstance3.delayedCh_BZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38589),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.delayedCh_A_2_LC_10_11_2 .C_ON=1'b0;
    defparam \QuadInstance3.delayedCh_A_2_LC_10_11_2 .SEQ_MODE=4'b1000;
    defparam \QuadInstance3.delayedCh_A_2_LC_10_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance3.delayedCh_A_2_LC_10_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19068),
            .lcout(\QuadInstance3.delayedCh_AZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38589),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.delayedCh_A_1_LC_10_11_3 .C_ON=1'b0;
    defparam \QuadInstance3.delayedCh_A_1_LC_10_11_3 .SEQ_MODE=4'b1000;
    defparam \QuadInstance3.delayedCh_A_1_LC_10_11_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \QuadInstance3.delayedCh_A_1_LC_10_11_3  (
            .in0(N__20388),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\QuadInstance3.delayedCh_AZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38589),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_RNIEUAL1_7_LC_10_11_4 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_RNIEUAL1_7_LC_10_11_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNIEUAL1_7_LC_10_11_4 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance3.Quad_RNIEUAL1_7_LC_10_11_4  (
            .in0(N__26336),
            .in1(N__21933),
            .in2(N__18975),
            .in3(N__19027),
            .lcout(\QuadInstance3.Quad_RNIEUAL1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.Quad_RNO_0_15_LC_10_11_5 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_RNO_0_15_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance3.Quad_RNO_0_15_LC_10_11_5 .LUT_INIT=16'b0011110010011100;
    LogicCell40 \QuadInstance3.Quad_RNO_0_15_LC_10_11_5  (
            .in0(N__19029),
            .in1(N__24335),
            .in2(N__18977),
            .in3(N__21935),
            .lcout(\QuadInstance3.un1_Quad_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam quadWrite_3_LC_10_11_6.C_ON=1'b0;
    defparam quadWrite_3_LC_10_11_6.SEQ_MODE=4'b1000;
    defparam quadWrite_3_LC_10_11_6.LUT_INIT=16'b0010000000000000;
    LogicCell40 quadWrite_3_LC_10_11_6 (
            .in0(N__23444),
            .in1(N__33822),
            .in2(N__33661),
            .in3(N__33436),
            .lcout(quadWriteZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38589),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance3.delayedCh_B_1_LC_10_11_7 .C_ON=1'b0;
    defparam \QuadInstance3.delayedCh_B_1_LC_10_11_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance3.delayedCh_B_1_LC_10_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance3.delayedCh_B_1_LC_10_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18879),
            .lcout(\QuadInstance3.delayedCh_BZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38589),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_10_12_0 .C_ON=1'b0;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_10_12_0 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance5.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_10_12_0  (
            .in0(N__19179),
            .in1(N__19198),
            .in2(N__19394),
            .in3(N__19185),
            .lcout(\PWMInstance5.un1_PWMPulseWidthCount_0_I_15_c_RNO_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.periodCounter_RNI5J7E_14_LC_10_12_1 .C_ON=1'b0;
    defparam \PWMInstance5.periodCounter_RNI5J7E_14_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance5.periodCounter_RNI5J7E_14_LC_10_12_1 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \PWMInstance5.periodCounter_RNI5J7E_14_LC_10_12_1  (
            .in0(N__19255),
            .in1(N__19237),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\PWMInstance5.un1_periodCounter12_1_0_a2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.periodCounter_RNIIJIT_10_LC_10_12_2 .C_ON=1'b0;
    defparam \PWMInstance5.periodCounter_RNIIJIT_10_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \PWMInstance5.periodCounter_RNIIJIT_10_LC_10_12_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \PWMInstance5.periodCounter_RNIIJIT_10_LC_10_12_2  (
            .in0(N__19172),
            .in1(N__19219),
            .in2(N__19203),
            .in3(N__19199),
            .lcout(\PWMInstance5.un1_periodCounter12_1_0_a2_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.PWMPulseWidthCount_esr_4_LC_10_12_3 .C_ON=1'b0;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_4_LC_10_12_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_4_LC_10_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance5.PWMPulseWidthCount_esr_4_LC_10_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36494),
            .lcout(\PWMInstance5.PWMPulseWidthCountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38578),
            .ce(N__19597),
            .sr(N__35739));
    defparam \PWMInstance5.PWMPulseWidthCount_esr_5_LC_10_12_4 .C_ON=1'b0;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_5_LC_10_12_4 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_5_LC_10_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance5.PWMPulseWidthCount_esr_5_LC_10_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36366),
            .lcout(\PWMInstance5.PWMPulseWidthCountZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38578),
            .ce(N__19597),
            .sr(N__35739));
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_10_12_5 .C_ON=1'b0;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_10_12_5 .SEQ_MODE=4'b0000;
    defparam \PWMInstance5.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_10_12_5 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance5.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_10_12_5  (
            .in0(N__19128),
            .in1(N__19171),
            .in2(N__19370),
            .in3(N__19158),
            .lcout(\PWMInstance5.un1_PWMPulseWidthCount_0_I_33_c_RNO_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.PWMPulseWidthCount_esr_11_LC_10_12_7 .C_ON=1'b0;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_11_LC_10_12_7 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_11_LC_10_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance5.PWMPulseWidthCount_esr_11_LC_10_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36004),
            .lcout(\PWMInstance5.PWMPulseWidthCountZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38578),
            .ce(N__19597),
            .sr(N__35739));
    defparam \PWMInstance5.out_RNO_0_LC_10_13_0 .C_ON=1'b0;
    defparam \PWMInstance5.out_RNO_0_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance5.out_RNO_0_LC_10_13_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \PWMInstance5.out_RNO_0_LC_10_13_0  (
            .in0(N__19570),
            .in1(N__19552),
            .in2(N__20244),
            .in3(N__19316),
            .lcout(\PWMInstance5.un1_periodCounter12_1_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.clkCount_0_LC_10_13_1 .C_ON=1'b0;
    defparam \PWMInstance5.clkCount_0_LC_10_13_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.clkCount_0_LC_10_13_1 .LUT_INIT=16'b1010000010100101;
    LogicCell40 \PWMInstance5.clkCount_0_LC_10_13_1  (
            .in0(N__19553),
            .in1(_gnd_net_),
            .in2(N__20231),
            .in3(N__19571),
            .lcout(\PWMInstance5.clkCountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38568),
            .ce(),
            .sr(N__35747));
    defparam \PWMInstance5.PWMPulseWidthCount_esr_ctle_15_LC_10_13_2 .C_ON=1'b0;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_ctle_15_LC_10_13_2 .SEQ_MODE=4'b0000;
    defparam \PWMInstance5.PWMPulseWidthCount_esr_ctle_15_LC_10_13_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \PWMInstance5.PWMPulseWidthCount_esr_ctle_15_LC_10_13_2  (
            .in0(_gnd_net_),
            .in1(N__35827),
            .in2(_gnd_net_),
            .in3(N__20224),
            .lcout(\PWMInstance5.pwmWrite_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.clkCount_1_LC_10_13_3 .C_ON=1'b0;
    defparam \PWMInstance5.clkCount_1_LC_10_13_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance5.clkCount_1_LC_10_13_3 .LUT_INIT=16'b1111000000001010;
    LogicCell40 \PWMInstance5.clkCount_1_LC_10_13_3  (
            .in0(N__19554),
            .in1(_gnd_net_),
            .in2(N__20232),
            .in3(N__19572),
            .lcout(\PWMInstance5.clkCountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38568),
            .ce(),
            .sr(N__35747));
    defparam \PWMInstance5.clkCount_RNI8JO8_0_LC_10_13_4 .C_ON=1'b0;
    defparam \PWMInstance5.clkCount_RNI8JO8_0_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance5.clkCount_RNI8JO8_0_LC_10_13_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \PWMInstance5.clkCount_RNI8JO8_0_LC_10_13_4  (
            .in0(N__20240),
            .in1(N__19569),
            .in2(_gnd_net_),
            .in3(N__19551),
            .lcout(\PWMInstance5.periodCounter12 ),
            .ltout(\PWMInstance5.periodCounter12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.periodCounter_RNIP0851_15_LC_10_13_5 .C_ON=1'b0;
    defparam \PWMInstance5.periodCounter_RNIP0851_15_LC_10_13_5 .SEQ_MODE=4'b0000;
    defparam \PWMInstance5.periodCounter_RNIP0851_15_LC_10_13_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \PWMInstance5.periodCounter_RNIP0851_15_LC_10_13_5  (
            .in0(N__19519),
            .in1(N__19501),
            .in2(N__19482),
            .in3(N__19278),
            .lcout(),
            .ltout(\PWMInstance5.un1_periodCounter12_1_0_a2_0_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.periodCounter_RNI8HQJ4_10_LC_10_13_6 .C_ON=1'b0;
    defparam \PWMInstance5.periodCounter_RNI8HQJ4_10_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \PWMInstance5.periodCounter_RNI8HQJ4_10_LC_10_13_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \PWMInstance5.periodCounter_RNI8HQJ4_10_LC_10_13_6  (
            .in0(N__19323),
            .in1(N__19479),
            .in2(N__19470),
            .in3(N__19467),
            .lcout(\PWMInstance5.out_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.periodCounter_RNIVUF81_11_LC_10_14_4 .C_ON=1'b0;
    defparam \PWMInstance5.periodCounter_RNIVUF81_11_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance5.periodCounter_RNIVUF81_11_LC_10_14_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \PWMInstance5.periodCounter_RNIVUF81_11_LC_10_14_4  (
            .in0(N__19414),
            .in1(N__19395),
            .in2(N__19371),
            .in3(N__19347),
            .lcout(\PWMInstance5.un1_periodCounter12_1_0_a2_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance5.periodCounter_RNICQ7E_16_LC_10_14_7 .C_ON=1'b0;
    defparam \PWMInstance5.periodCounter_RNICQ7E_16_LC_10_14_7 .SEQ_MODE=4'b0000;
    defparam \PWMInstance5.periodCounter_RNICQ7E_16_LC_10_14_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \PWMInstance5.periodCounter_RNICQ7E_16_LC_10_14_7  (
            .in0(_gnd_net_),
            .in1(N__19315),
            .in2(_gnd_net_),
            .in3(N__19299),
            .lcout(\PWMInstance5.un1_periodCounter12_1_0_a2_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance6.periodCounter_RNI7M9F_14_LC_10_15_0 .C_ON=1'b0;
    defparam \PWMInstance6.periodCounter_RNI7M9F_14_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance6.periodCounter_RNI7M9F_14_LC_10_15_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \PWMInstance6.periodCounter_RNI7M9F_14_LC_10_15_0  (
            .in0(N__23167),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20210),
            .lcout(),
            .ltout(\PWMInstance6.un1_periodCounter12_1_0_a2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance6.periodCounter_RNINBG41_10_LC_10_15_1 .C_ON=1'b0;
    defparam \PWMInstance6.periodCounter_RNINBG41_10_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance6.periodCounter_RNINBG41_10_LC_10_15_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \PWMInstance6.periodCounter_RNINBG41_10_LC_10_15_1  (
            .in0(N__23053),
            .in1(N__23128),
            .in2(N__19710),
            .in3(N__20351),
            .lcout(),
            .ltout(\PWMInstance6.un1_periodCounter12_1_0_a2_0_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance6.periodCounter_RNISI7C4_10_LC_10_15_2 .C_ON=1'b0;
    defparam \PWMInstance6.periodCounter_RNISI7C4_10_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \PWMInstance6.periodCounter_RNISI7C4_10_LC_10_15_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \PWMInstance6.periodCounter_RNISI7C4_10_LC_10_15_2  (
            .in0(N__19704),
            .in1(N__21099),
            .in2(N__19707),
            .in3(N__21138),
            .lcout(\PWMInstance6.out_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance6.periodCounter_RNI34321_11_LC_10_15_4 .C_ON=1'b0;
    defparam \PWMInstance6.periodCounter_RNI34321_11_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance6.periodCounter_RNI34321_11_LC_10_15_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \PWMInstance6.periodCounter_RNI34321_11_LC_10_15_4  (
            .in0(N__21226),
            .in1(N__20323),
            .in2(N__23102),
            .in3(N__20179),
            .lcout(\PWMInstance6.un1_periodCounter12_1_0_a2_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_10_16_1 .C_ON=1'b0;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_10_16_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_10_16_1 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance6.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_10_16_1  (
            .in0(N__19692),
            .in1(N__19698),
            .in2(N__20187),
            .in3(N__20211),
            .lcout(\PWMInstance6.un1_PWMPulseWidthCount_0_I_9_c_RNO_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance6.PWMPulseWidthCount_esr_2_LC_10_16_2 .C_ON=1'b0;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_2_LC_10_16_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_2_LC_10_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance6.PWMPulseWidthCount_esr_2_LC_10_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31592),
            .lcout(\PWMInstance6.PWMPulseWidthCountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38550),
            .ce(N__24556),
            .sr(N__35763));
    defparam \PWMInstance6.PWMPulseWidthCount_esr_3_LC_10_16_3 .C_ON=1'b0;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_3_LC_10_16_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_3_LC_10_16_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \PWMInstance6.PWMPulseWidthCount_esr_3_LC_10_16_3  (
            .in0(_gnd_net_),
            .in1(N__32072),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PWMInstance6.PWMPulseWidthCountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38550),
            .ce(N__24556),
            .sr(N__35763));
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_10_16_6 .C_ON=1'b0;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_10_16_6 .SEQ_MODE=4'b0000;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_10_16_6 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance6.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_10_16_6  (
            .in0(N__20355),
            .in1(N__22959),
            .in2(N__19686),
            .in3(N__20328),
            .lcout(\PWMInstance6.un1_PWMPulseWidthCount_0_I_15_c_RNO_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance6.PWMPulseWidthCount_esr_4_LC_10_16_7 .C_ON=1'b0;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_4_LC_10_16_7 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_4_LC_10_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance6.PWMPulseWidthCount_esr_4_LC_10_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36512),
            .lcout(\PWMInstance6.PWMPulseWidthCountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38550),
            .ce(N__24556),
            .sr(N__35763));
    defparam \QuadInstance2.Quad_2_LC_11_4_1 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_2_LC_11_4_1 .SEQ_MODE=4'b1000;
    defparam \QuadInstance2.Quad_2_LC_11_4_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance2.Quad_2_LC_11_4_1  (
            .in0(N__31587),
            .in1(N__22192),
            .in2(_gnd_net_),
            .in3(N__19677),
            .lcout(dataRead2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38673),
            .ce(),
            .sr(N__35690));
    defparam \QuadInstance3.Quad_2_LC_11_4_2 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_2_LC_11_4_2 .SEQ_MODE=4'b1000;
    defparam \QuadInstance3.Quad_2_LC_11_4_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance3.Quad_2_LC_11_4_2  (
            .in0(N__31589),
            .in1(N__22019),
            .in2(_gnd_net_),
            .in3(N__19665),
            .lcout(dataRead3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38673),
            .ce(),
            .sr(N__35690));
    defparam \QuadInstance2.Quad_6_LC_11_4_3 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_6_LC_11_4_3 .SEQ_MODE=4'b1000;
    defparam \QuadInstance2.Quad_6_LC_11_4_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance2.Quad_6_LC_11_4_3  (
            .in0(N__31120),
            .in1(N__22194),
            .in2(_gnd_net_),
            .in3(N__19770),
            .lcout(dataRead2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38673),
            .ce(),
            .sr(N__35690));
    defparam \QuadInstance6.Quad_2_LC_11_4_4 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_2_LC_11_4_4 .SEQ_MODE=4'b1000;
    defparam \QuadInstance6.Quad_2_LC_11_4_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance6.Quad_2_LC_11_4_4  (
            .in0(N__31590),
            .in1(N__22798),
            .in2(_gnd_net_),
            .in3(N__20430),
            .lcout(dataRead6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38673),
            .ce(),
            .sr(N__35690));
    defparam \QuadInstance7.Quad_2_LC_11_4_5 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_2_LC_11_4_5 .SEQ_MODE=4'b1000;
    defparam \QuadInstance7.Quad_2_LC_11_4_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance7.Quad_2_LC_11_4_5  (
            .in0(N__31588),
            .in1(N__26052),
            .in2(_gnd_net_),
            .in3(N__19758),
            .lcout(dataRead7_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38673),
            .ce(),
            .sr(N__35690));
    defparam \QuadInstance1.Quad_3_LC_11_4_6 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_3_LC_11_4_6 .SEQ_MODE=4'b1000;
    defparam \QuadInstance1.Quad_3_LC_11_4_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance1.Quad_3_LC_11_4_6  (
            .in0(N__24098),
            .in1(N__32086),
            .in2(_gnd_net_),
            .in3(N__21615),
            .lcout(dataRead1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38673),
            .ce(),
            .sr(N__35690));
    defparam \QuadInstance2.Quad_3_LC_11_4_7 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_3_LC_11_4_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance2.Quad_3_LC_11_4_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance2.Quad_3_LC_11_4_7  (
            .in0(N__32087),
            .in1(N__22193),
            .in2(_gnd_net_),
            .in3(N__19746),
            .lcout(dataRead2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38673),
            .ce(),
            .sr(N__35690));
    defparam \QuadInstance5.Quad_4_LC_11_5_0 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_4_LC_11_5_0 .SEQ_MODE=4'b1000;
    defparam \QuadInstance5.Quad_4_LC_11_5_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance5.Quad_4_LC_11_5_0  (
            .in0(N__36514),
            .in1(N__25800),
            .in2(_gnd_net_),
            .in3(N__19734),
            .lcout(dataRead5_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38662),
            .ce(),
            .sr(N__35692));
    defparam \QuadInstance5.Quad_6_LC_11_5_1 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_6_LC_11_5_1 .SEQ_MODE=4'b1000;
    defparam \QuadInstance5.Quad_6_LC_11_5_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance5.Quad_6_LC_11_5_1  (
            .in0(N__25798),
            .in1(N__31112),
            .in2(_gnd_net_),
            .in3(N__19728),
            .lcout(dataRead5_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38662),
            .ce(),
            .sr(N__35692));
    defparam \QuadInstance6.Quad_6_LC_11_5_2 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_6_LC_11_5_2 .SEQ_MODE=4'b1000;
    defparam \QuadInstance6.Quad_6_LC_11_5_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance6.Quad_6_LC_11_5_2  (
            .in0(N__31113),
            .in1(N__22796),
            .in2(_gnd_net_),
            .in3(N__20508),
            .lcout(dataRead6_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38662),
            .ce(),
            .sr(N__35692));
    defparam \QuadInstance7.Quad_6_LC_11_5_3 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_6_LC_11_5_3 .SEQ_MODE=4'b1000;
    defparam \QuadInstance7.Quad_6_LC_11_5_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance7.Quad_6_LC_11_5_3  (
            .in0(N__31110),
            .in1(N__26014),
            .in2(_gnd_net_),
            .in3(N__19722),
            .lcout(dataRead7_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38662),
            .ce(),
            .sr(N__35692));
    defparam \QuadInstance7.Quad_9_LC_11_5_4 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_9_LC_11_5_4 .SEQ_MODE=4'b1000;
    defparam \QuadInstance7.Quad_9_LC_11_5_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance7.Quad_9_LC_11_5_4  (
            .in0(N__26013),
            .in1(N__28572),
            .in2(_gnd_net_),
            .in3(N__19836),
            .lcout(dataRead7_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38662),
            .ce(),
            .sr(N__35692));
    defparam \QuadInstance5.Quad_8_LC_11_5_5 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_8_LC_11_5_5 .SEQ_MODE=4'b1000;
    defparam \QuadInstance5.Quad_8_LC_11_5_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance5.Quad_8_LC_11_5_5  (
            .in0(N__25799),
            .in1(N__28988),
            .in2(_gnd_net_),
            .in3(N__19824),
            .lcout(dataRead5_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38662),
            .ce(),
            .sr(N__35692));
    defparam \QuadInstance6.Quad_8_LC_11_5_6 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_8_LC_11_5_6 .SEQ_MODE=4'b1000;
    defparam \QuadInstance6.Quad_8_LC_11_5_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance6.Quad_8_LC_11_5_6  (
            .in0(N__28989),
            .in1(N__22797),
            .in2(_gnd_net_),
            .in3(N__20490),
            .lcout(dataRead6_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38662),
            .ce(),
            .sr(N__35692));
    defparam \QuadInstance3.Quad_3_LC_11_5_7 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_3_LC_11_5_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance3.Quad_3_LC_11_5_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance3.Quad_3_LC_11_5_7  (
            .in0(N__32073),
            .in1(N__22018),
            .in2(_gnd_net_),
            .in3(N__19815),
            .lcout(dataRead3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38662),
            .ce(),
            .sr(N__35692));
    defparam \QuadInstance1.Quad_7_LC_11_6_0 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_7_LC_11_6_0 .SEQ_MODE=4'b1000;
    defparam \QuadInstance1.Quad_7_LC_11_6_0 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \QuadInstance1.Quad_7_LC_11_6_0  (
            .in0(N__29448),
            .in1(_gnd_net_),
            .in2(N__24099),
            .in3(N__21564),
            .lcout(dataRead1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38650),
            .ce(),
            .sr(N__35700));
    defparam \QuadInstance2.Quad_7_LC_11_6_1 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_7_LC_11_6_1 .SEQ_MODE=4'b1000;
    defparam \QuadInstance2.Quad_7_LC_11_6_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance2.Quad_7_LC_11_6_1  (
            .in0(N__29449),
            .in1(N__22185),
            .in2(_gnd_net_),
            .in3(N__19803),
            .lcout(dataRead2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38650),
            .ce(),
            .sr(N__35700));
    defparam \QuadInstance3.Quad_7_LC_11_6_2 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_7_LC_11_6_2 .SEQ_MODE=4'b1000;
    defparam \QuadInstance3.Quad_7_LC_11_6_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance3.Quad_7_LC_11_6_2  (
            .in0(N__22015),
            .in1(N__29450),
            .in2(_gnd_net_),
            .in3(N__19794),
            .lcout(dataRead3_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38650),
            .ce(),
            .sr(N__35700));
    defparam \QuadInstance5.Quad_7_LC_11_6_3 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_7_LC_11_6_3 .SEQ_MODE=4'b1000;
    defparam \QuadInstance5.Quad_7_LC_11_6_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance5.Quad_7_LC_11_6_3  (
            .in0(N__29451),
            .in1(N__25772),
            .in2(_gnd_net_),
            .in3(N__19785),
            .lcout(dataRead5_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38650),
            .ce(),
            .sr(N__35700));
    defparam \QuadInstance3.Quad_5_LC_11_6_4 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_5_LC_11_6_4 .SEQ_MODE=4'b1000;
    defparam \QuadInstance3.Quad_5_LC_11_6_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance3.Quad_5_LC_11_6_4  (
            .in0(N__22014),
            .in1(N__36368),
            .in2(_gnd_net_),
            .in3(N__19779),
            .lcout(dataRead3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38650),
            .ce(),
            .sr(N__35700));
    defparam \QuadInstance7.Quad_7_LC_11_6_5 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_7_LC_11_6_5 .SEQ_MODE=4'b1000;
    defparam \QuadInstance7.Quad_7_LC_11_6_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance7.Quad_7_LC_11_6_5  (
            .in0(N__29452),
            .in1(N__26012),
            .in2(_gnd_net_),
            .in3(N__19890),
            .lcout(dataRead7_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38650),
            .ce(),
            .sr(N__35700));
    defparam \QuadInstance1.Quad_8_LC_11_6_6 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_8_LC_11_6_6 .SEQ_MODE=4'b1000;
    defparam \QuadInstance1.Quad_8_LC_11_6_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance1.Quad_8_LC_11_6_6  (
            .in0(N__24080),
            .in1(N__28987),
            .in2(_gnd_net_),
            .in3(N__21552),
            .lcout(dataRead1_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38650),
            .ce(),
            .sr(N__35700));
    defparam \QuadInstance6.Quad_11_LC_11_6_7 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_11_LC_11_6_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance6.Quad_11_LC_11_6_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \QuadInstance6.Quad_11_LC_11_6_7  (
            .in0(N__35993),
            .in1(_gnd_net_),
            .in2(N__22805),
            .in3(N__20475),
            .lcout(dataRead6_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38650),
            .ce(),
            .sr(N__35700));
    defparam \QuadInstance0.Quad_11_LC_11_7_0 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_11_LC_11_7_0 .SEQ_MODE=4'b1000;
    defparam \QuadInstance0.Quad_11_LC_11_7_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance0.Quad_11_LC_11_7_0  (
            .in0(N__36005),
            .in1(N__33132),
            .in2(_gnd_net_),
            .in3(N__30066),
            .lcout(dataRead0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38641),
            .ce(),
            .sr(N__35705));
    defparam \QuadInstance1.Quad_11_LC_11_7_1 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_11_LC_11_7_1 .SEQ_MODE=4'b1000;
    defparam \QuadInstance1.Quad_11_LC_11_7_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance1.Quad_11_LC_11_7_1  (
            .in0(N__24095),
            .in1(N__36006),
            .in2(_gnd_net_),
            .in3(N__21675),
            .lcout(dataRead1_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38641),
            .ce(),
            .sr(N__35705));
    defparam \QuadInstance2.Quad_11_LC_11_7_2 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_11_LC_11_7_2 .SEQ_MODE=4'b1000;
    defparam \QuadInstance2.Quad_11_LC_11_7_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \QuadInstance2.Quad_11_LC_11_7_2  (
            .in0(N__22186),
            .in1(_gnd_net_),
            .in2(N__36015),
            .in3(N__19878),
            .lcout(dataRead2_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38641),
            .ce(),
            .sr(N__35705));
    defparam \QuadInstance5.Quad_10_LC_11_7_3 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_10_LC_11_7_3 .SEQ_MODE=4'b1000;
    defparam \QuadInstance5.Quad_10_LC_11_7_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance5.Quad_10_LC_11_7_3  (
            .in0(N__25796),
            .in1(N__36142),
            .in2(_gnd_net_),
            .in3(N__19869),
            .lcout(dataRead5_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38641),
            .ce(),
            .sr(N__35705));
    defparam \QuadInstance5.Quad_11_LC_11_7_4 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_11_LC_11_7_4 .SEQ_MODE=4'b1000;
    defparam \QuadInstance5.Quad_11_LC_11_7_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance5.Quad_11_LC_11_7_4  (
            .in0(N__36010),
            .in1(N__25797),
            .in2(_gnd_net_),
            .in3(N__19863),
            .lcout(dataRead5_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38641),
            .ce(),
            .sr(N__35705));
    defparam \QuadInstance2.Quad_8_LC_11_7_5 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_8_LC_11_7_5 .SEQ_MODE=4'b1000;
    defparam \QuadInstance2.Quad_8_LC_11_7_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance2.Quad_8_LC_11_7_5  (
            .in0(N__28986),
            .in1(N__22187),
            .in2(_gnd_net_),
            .in3(N__19857),
            .lcout(dataRead2_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38641),
            .ce(),
            .sr(N__35705));
    defparam \QuadInstance3.Quad_9_LC_11_7_6 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_9_LC_11_7_6 .SEQ_MODE=4'b1000;
    defparam \QuadInstance3.Quad_9_LC_11_7_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance3.Quad_9_LC_11_7_6  (
            .in0(N__28559),
            .in1(N__22017),
            .in2(_gnd_net_),
            .in3(N__19845),
            .lcout(dataRead3_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38641),
            .ce(),
            .sr(N__35705));
    defparam \QuadInstance0.Quad_3_LC_11_7_7 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_3_LC_11_7_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance0.Quad_3_LC_11_7_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance0.Quad_3_LC_11_7_7  (
            .in0(N__33131),
            .in1(N__32050),
            .in2(_gnd_net_),
            .in3(N__29865),
            .lcout(dataRead0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38641),
            .ce(),
            .sr(N__35705));
    defparam OutReg_ess_RNO_3_13_LC_11_8_2.C_ON=1'b0;
    defparam OutReg_ess_RNO_3_13_LC_11_8_2.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_3_13_LC_11_8_2.LUT_INIT=16'b0101001001010111;
    LogicCell40 OutReg_ess_RNO_3_13_LC_11_8_2 (
            .in0(N__28013),
            .in1(N__19921),
            .in2(N__28133),
            .in3(N__19960),
            .lcout(OutReg_0_4_i_m3_ns_1_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_2_13_LC_11_8_3.C_ON=1'b0;
    defparam OutReg_ess_RNO_2_13_LC_11_8_3.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_2_13_LC_11_8_3.LUT_INIT=16'b1000100011110011;
    LogicCell40 OutReg_ess_RNO_2_13_LC_11_8_3 (
            .in0(N__23922),
            .in1(N__38152),
            .in2(N__20019),
            .in3(N__27543),
            .lcout(OutReg_ess_RNO_2Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.Quad_13_LC_11_8_4 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_13_LC_11_8_4 .SEQ_MODE=4'b1000;
    defparam \QuadInstance2.Quad_13_LC_11_8_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance2.Quad_13_LC_11_8_4  (
            .in0(N__28684),
            .in1(N__22188),
            .in2(_gnd_net_),
            .in3(N__19986),
            .lcout(dataRead2_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38631),
            .ce(),
            .sr(N__35714));
    defparam \QuadInstance3.Quad_13_LC_11_8_5 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_13_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \QuadInstance3.Quad_13_LC_11_8_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance3.Quad_13_LC_11_8_5  (
            .in0(N__22016),
            .in1(N__28685),
            .in2(_gnd_net_),
            .in3(N__19944),
            .lcout(dataRead3_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38631),
            .ce(),
            .sr(N__35714));
    defparam \QuadInstance6.Quad_13_LC_11_8_6 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_13_LC_11_8_6 .SEQ_MODE=4'b1000;
    defparam \QuadInstance6.Quad_13_LC_11_8_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance6.Quad_13_LC_11_8_6  (
            .in0(N__28686),
            .in1(N__22755),
            .in2(_gnd_net_),
            .in3(N__20625),
            .lcout(dataRead6_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38631),
            .ce(),
            .sr(N__35714));
    defparam \QuadInstance3.Quad_12_LC_11_9_0 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_12_LC_11_9_0 .SEQ_MODE=4'b1000;
    defparam \QuadInstance3.Quad_12_LC_11_9_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance3.Quad_12_LC_11_9_0  (
            .in0(N__28800),
            .in1(N__22003),
            .in2(_gnd_net_),
            .in3(N__19905),
            .lcout(dataRead3_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38618),
            .ce(),
            .sr(N__35721));
    defparam \QuadInstance6.Quad_12_LC_11_9_1 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_12_LC_11_9_1 .SEQ_MODE=4'b1000;
    defparam \QuadInstance6.Quad_12_LC_11_9_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance6.Quad_12_LC_11_9_1  (
            .in0(N__28801),
            .in1(N__22754),
            .in2(_gnd_net_),
            .in3(N__20466),
            .lcout(dataRead6_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38618),
            .ce(),
            .sr(N__35721));
    defparam \QuadInstance3.Quad_8_LC_11_9_2 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_8_LC_11_9_2 .SEQ_MODE=4'b1000;
    defparam \QuadInstance3.Quad_8_LC_11_9_2 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \QuadInstance3.Quad_8_LC_11_9_2  (
            .in0(N__28952),
            .in1(_gnd_net_),
            .in2(N__19899),
            .in3(N__22004),
            .lcout(dataRead3_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38618),
            .ce(),
            .sr(N__35721));
    defparam \QuadInstance3.Quad_14_LC_11_9_3 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_14_LC_11_9_3 .SEQ_MODE=4'b1000;
    defparam \QuadInstance3.Quad_14_LC_11_9_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance3.Quad_14_LC_11_9_3  (
            .in0(N__22000),
            .in1(N__34365),
            .in2(_gnd_net_),
            .in3(N__20157),
            .lcout(dataRead3_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38618),
            .ce(),
            .sr(N__35721));
    defparam \QuadInstance5.Quad_2_LC_11_9_4 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_2_LC_11_9_4 .SEQ_MODE=4'b1000;
    defparam \QuadInstance5.Quad_2_LC_11_9_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance5.Quad_2_LC_11_9_4  (
            .in0(N__31542),
            .in1(N__25806),
            .in2(_gnd_net_),
            .in3(N__20151),
            .lcout(dataRead5_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38618),
            .ce(),
            .sr(N__35721));
    defparam \QuadInstance7.Quad_14_LC_11_9_5 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_14_LC_11_9_5 .SEQ_MODE=4'b1000;
    defparam \QuadInstance7.Quad_14_LC_11_9_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance7.Quad_14_LC_11_9_5  (
            .in0(N__34366),
            .in1(N__26038),
            .in2(_gnd_net_),
            .in3(N__20142),
            .lcout(dataRead7_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38618),
            .ce(),
            .sr(N__35721));
    defparam \QuadInstance3.Quad_10_LC_11_9_6 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_10_LC_11_9_6 .SEQ_MODE=4'b1000;
    defparam \QuadInstance3.Quad_10_LC_11_9_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance3.Quad_10_LC_11_9_6  (
            .in0(N__36089),
            .in1(N__22002),
            .in2(_gnd_net_),
            .in3(N__20133),
            .lcout(dataRead3_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38618),
            .ce(),
            .sr(N__35721));
    defparam \QuadInstance3.Quad_11_LC_11_9_7 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_11_LC_11_9_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance3.Quad_11_LC_11_9_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \QuadInstance3.Quad_11_LC_11_9_7  (
            .in0(N__22001),
            .in1(_gnd_net_),
            .in2(N__35973),
            .in3(N__20127),
            .lcout(dataRead3_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38618),
            .ce(),
            .sr(N__35721));
    defparam OutReg_ess_RNO_0_13_LC_11_10_0.C_ON=1'b0;
    defparam OutReg_ess_RNO_0_13_LC_11_10_0.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_0_13_LC_11_10_0.LUT_INIT=16'b1110111001000100;
    LogicCell40 OutReg_ess_RNO_0_13_LC_11_10_0 (
            .in0(N__37558),
            .in1(N__20121),
            .in2(_gnd_net_),
            .in3(N__20730),
            .lcout(OutReg_ess_RNO_0Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_4_11_LC_11_10_1.C_ON=1'b0;
    defparam OutReg_ess_RNO_4_11_LC_11_10_1.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_4_11_LC_11_10_1.LUT_INIT=16'b0000010110111011;
    LogicCell40 OutReg_ess_RNO_4_11_LC_11_10_1 (
            .in0(N__28015),
            .in1(N__30097),
            .in2(N__25122),
            .in3(N__28137),
            .lcout(),
            .ltout(OutReg_0_5_i_m3_i_m3_ns_1_11_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_2_11_LC_11_10_2.C_ON=1'b0;
    defparam OutReg_ess_RNO_2_11_LC_11_10_2.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_2_11_LC_11_10_2.LUT_INIT=16'b1100101100001011;
    LogicCell40 OutReg_ess_RNO_2_11_LC_11_10_2 (
            .in0(N__20108),
            .in1(N__32948),
            .in2(N__20082),
            .in3(N__23366),
            .lcout(OutReg_ess_RNO_2Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_esr_RNO_3_14_LC_11_10_4.C_ON=1'b0;
    defparam OutReg_esr_RNO_3_14_LC_11_10_4.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_3_14_LC_11_10_4.LUT_INIT=16'b0000010111110011;
    LogicCell40 OutReg_esr_RNO_3_14_LC_11_10_4 (
            .in0(N__20065),
            .in1(N__20048),
            .in2(N__28140),
            .in3(N__28014),
            .lcout(),
            .ltout(OutReg_0_4_i_m3_ns_1_14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_esr_RNO_1_14_LC_11_10_5.C_ON=1'b0;
    defparam OutReg_esr_RNO_1_14_LC_11_10_5.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_1_14_LC_11_10_5.LUT_INIT=16'b1100101000001111;
    LogicCell40 OutReg_esr_RNO_1_14_LC_11_10_5 (
            .in0(N__20263),
            .in1(N__20558),
            .in2(N__20247),
            .in3(N__37741),
            .lcout(OutReg_esr_RNO_1Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwmWrite_4_LC_11_11_4.C_ON=1'b0;
    defparam pwmWrite_4_LC_11_11_4.SEQ_MODE=4'b1000;
    defparam pwmWrite_4_LC_11_11_4.LUT_INIT=16'b0000001000000000;
    LogicCell40 pwmWrite_4_LC_11_11_4 (
            .in0(N__33749),
            .in1(N__33560),
            .in2(N__33464),
            .in3(N__33207),
            .lcout(pwmWriteZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38597),
            .ce(),
            .sr(_gnd_net_));
    defparam data_received_esr_4_LC_11_12_3.C_ON=1'b0;
    defparam data_received_esr_4_LC_11_12_3.SEQ_MODE=4'b1000;
    defparam data_received_esr_4_LC_11_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 data_received_esr_4_LC_11_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30621),
            .lcout(data_receivedZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38590),
            .ce(N__26184),
            .sr(N__26154));
    defparam pwmWrite_fast_5_LC_11_13_4.C_ON=1'b0;
    defparam pwmWrite_fast_5_LC_11_13_4.SEQ_MODE=4'b1000;
    defparam pwmWrite_fast_5_LC_11_13_4.LUT_INIT=16'b0000001000000000;
    LogicCell40 pwmWrite_fast_5_LC_11_13_4 (
            .in0(N__23429),
            .in1(N__33440),
            .in2(N__33600),
            .in3(N__33751),
            .lcout(pwmWrite_fastZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38579),
            .ce(),
            .sr(_gnd_net_));
    defparam pwmWrite_5_LC_11_13_5.C_ON=1'b0;
    defparam pwmWrite_5_LC_11_13_5.SEQ_MODE=4'b1000;
    defparam pwmWrite_5_LC_11_13_5.LUT_INIT=16'b0000001000000000;
    LogicCell40 pwmWrite_5_LC_11_13_5 (
            .in0(N__33750),
            .in1(N__33561),
            .in2(N__33465),
            .in3(N__23428),
            .lcout(pwmWriteZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38579),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance6.periodCounter_0_LC_11_14_0 .C_ON=1'b1;
    defparam \PWMInstance6.periodCounter_0_LC_11_14_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.periodCounter_0_LC_11_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance6.periodCounter_0_LC_11_14_0  (
            .in0(_gnd_net_),
            .in1(N__21090),
            .in2(N__21162),
            .in3(N__21158),
            .lcout(\PWMInstance6.periodCounterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_11_14_0_),
            .carryout(\PWMInstance6.un1_periodCounter_2_cry_0 ),
            .clk(N__38569),
            .ce(),
            .sr(N__35298));
    defparam \PWMInstance6.periodCounter_1_LC_11_14_1 .C_ON=1'b1;
    defparam \PWMInstance6.periodCounter_1_LC_11_14_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.periodCounter_1_LC_11_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance6.periodCounter_1_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(N__21074),
            .in2(_gnd_net_),
            .in3(N__20214),
            .lcout(\PWMInstance6.periodCounterZ0Z_1 ),
            .ltout(),
            .carryin(\PWMInstance6.un1_periodCounter_2_cry_0 ),
            .carryout(\PWMInstance6.un1_periodCounter_2_cry_1 ),
            .clk(N__38569),
            .ce(),
            .sr(N__35298));
    defparam \PWMInstance6.periodCounter_2_LC_11_14_2 .C_ON=1'b1;
    defparam \PWMInstance6.periodCounter_2_LC_11_14_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.periodCounter_2_LC_11_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance6.periodCounter_2_LC_11_14_2  (
            .in0(_gnd_net_),
            .in1(N__20209),
            .in2(_gnd_net_),
            .in3(N__20190),
            .lcout(\PWMInstance6.periodCounterZ0Z_2 ),
            .ltout(),
            .carryin(\PWMInstance6.un1_periodCounter_2_cry_1 ),
            .carryout(\PWMInstance6.un1_periodCounter_2_cry_2 ),
            .clk(N__38569),
            .ce(),
            .sr(N__35298));
    defparam \PWMInstance6.periodCounter_3_LC_11_14_3 .C_ON=1'b1;
    defparam \PWMInstance6.periodCounter_3_LC_11_14_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.periodCounter_3_LC_11_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance6.periodCounter_3_LC_11_14_3  (
            .in0(_gnd_net_),
            .in1(N__20180),
            .in2(_gnd_net_),
            .in3(N__20160),
            .lcout(\PWMInstance6.periodCounterZ0Z_3 ),
            .ltout(),
            .carryin(\PWMInstance6.un1_periodCounter_2_cry_2 ),
            .carryout(\PWMInstance6.un1_periodCounter_2_cry_3 ),
            .clk(N__38569),
            .ce(),
            .sr(N__35298));
    defparam \PWMInstance6.periodCounter_4_LC_11_14_4 .C_ON=1'b1;
    defparam \PWMInstance6.periodCounter_4_LC_11_14_4 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.periodCounter_4_LC_11_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance6.periodCounter_4_LC_11_14_4  (
            .in0(_gnd_net_),
            .in1(N__20350),
            .in2(_gnd_net_),
            .in3(N__20331),
            .lcout(\PWMInstance6.periodCounterZ0Z_4 ),
            .ltout(),
            .carryin(\PWMInstance6.un1_periodCounter_2_cry_3 ),
            .carryout(\PWMInstance6.un1_periodCounter_2_cry_4 ),
            .clk(N__38569),
            .ce(),
            .sr(N__35298));
    defparam \PWMInstance6.periodCounter_5_LC_11_14_5 .C_ON=1'b1;
    defparam \PWMInstance6.periodCounter_5_LC_11_14_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.periodCounter_5_LC_11_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance6.periodCounter_5_LC_11_14_5  (
            .in0(_gnd_net_),
            .in1(N__20327),
            .in2(_gnd_net_),
            .in3(N__20307),
            .lcout(\PWMInstance6.periodCounterZ0Z_5 ),
            .ltout(),
            .carryin(\PWMInstance6.un1_periodCounter_2_cry_4 ),
            .carryout(\PWMInstance6.un1_periodCounter_2_cry_5 ),
            .clk(N__38569),
            .ce(),
            .sr(N__35298));
    defparam \PWMInstance6.periodCounter_6_LC_11_14_6 .C_ON=1'b1;
    defparam \PWMInstance6.periodCounter_6_LC_11_14_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.periodCounter_6_LC_11_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance6.periodCounter_6_LC_11_14_6  (
            .in0(_gnd_net_),
            .in1(N__21041),
            .in2(_gnd_net_),
            .in3(N__20304),
            .lcout(\PWMInstance6.periodCounterZ0Z_6 ),
            .ltout(),
            .carryin(\PWMInstance6.un1_periodCounter_2_cry_5 ),
            .carryout(\PWMInstance6.un1_periodCounter_2_cry_6 ),
            .clk(N__38569),
            .ce(),
            .sr(N__35298));
    defparam \PWMInstance6.periodCounter_7_LC_11_14_7 .C_ON=1'b1;
    defparam \PWMInstance6.periodCounter_7_LC_11_14_7 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.periodCounter_7_LC_11_14_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance6.periodCounter_7_LC_11_14_7  (
            .in0(N__21422),
            .in1(N__21024),
            .in2(_gnd_net_),
            .in3(N__20301),
            .lcout(\PWMInstance6.periodCounterZ0Z_7 ),
            .ltout(),
            .carryin(\PWMInstance6.un1_periodCounter_2_cry_6 ),
            .carryout(\PWMInstance6.un1_periodCounter_2_cry_7 ),
            .clk(N__38569),
            .ce(),
            .sr(N__35298));
    defparam \PWMInstance6.periodCounter_8_LC_11_15_0 .C_ON=1'b1;
    defparam \PWMInstance6.periodCounter_8_LC_11_15_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.periodCounter_8_LC_11_15_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance6.periodCounter_8_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__21246),
            .in2(_gnd_net_),
            .in3(N__20298),
            .lcout(\PWMInstance6.periodCounterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_11_15_0_),
            .carryout(\PWMInstance6.un1_periodCounter_2_cry_8 ),
            .clk(N__38562),
            .ce(),
            .sr(N__35296));
    defparam \PWMInstance6.periodCounter_9_LC_11_15_1 .C_ON=1'b1;
    defparam \PWMInstance6.periodCounter_9_LC_11_15_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.periodCounter_9_LC_11_15_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance6.periodCounter_9_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(N__21227),
            .in2(_gnd_net_),
            .in3(N__20295),
            .lcout(\PWMInstance6.periodCounterZ0Z_9 ),
            .ltout(),
            .carryin(\PWMInstance6.un1_periodCounter_2_cry_8 ),
            .carryout(\PWMInstance6.un1_periodCounter_2_cry_9 ),
            .clk(N__38562),
            .ce(),
            .sr(N__35296));
    defparam \PWMInstance6.periodCounter_10_LC_11_15_2 .C_ON=1'b1;
    defparam \PWMInstance6.periodCounter_10_LC_11_15_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.periodCounter_10_LC_11_15_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance6.periodCounter_10_LC_11_15_2  (
            .in0(_gnd_net_),
            .in1(N__23129),
            .in2(_gnd_net_),
            .in3(N__20292),
            .lcout(\PWMInstance6.periodCounterZ0Z_10 ),
            .ltout(),
            .carryin(\PWMInstance6.un1_periodCounter_2_cry_9 ),
            .carryout(\PWMInstance6.un1_periodCounter_2_cry_10 ),
            .clk(N__38562),
            .ce(),
            .sr(N__35296));
    defparam \PWMInstance6.periodCounter_11_LC_11_15_3 .C_ON=1'b1;
    defparam \PWMInstance6.periodCounter_11_LC_11_15_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.periodCounter_11_LC_11_15_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance6.periodCounter_11_LC_11_15_3  (
            .in0(N__21420),
            .in1(N__23098),
            .in2(_gnd_net_),
            .in3(N__20289),
            .lcout(\PWMInstance6.periodCounterZ0Z_11 ),
            .ltout(),
            .carryin(\PWMInstance6.un1_periodCounter_2_cry_10 ),
            .carryout(\PWMInstance6.un1_periodCounter_2_cry_11 ),
            .clk(N__38562),
            .ce(),
            .sr(N__35296));
    defparam \PWMInstance6.periodCounter_12_LC_11_15_4 .C_ON=1'b1;
    defparam \PWMInstance6.periodCounter_12_LC_11_15_4 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.periodCounter_12_LC_11_15_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance6.periodCounter_12_LC_11_15_4  (
            .in0(N__21412),
            .in1(N__23054),
            .in2(_gnd_net_),
            .in3(N__20286),
            .lcout(\PWMInstance6.periodCounterZ0Z_12 ),
            .ltout(),
            .carryin(\PWMInstance6.un1_periodCounter_2_cry_11 ),
            .carryout(\PWMInstance6.un1_periodCounter_2_cry_12 ),
            .clk(N__38562),
            .ce(),
            .sr(N__35296));
    defparam \PWMInstance6.periodCounter_13_LC_11_15_5 .C_ON=1'b1;
    defparam \PWMInstance6.periodCounter_13_LC_11_15_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.periodCounter_13_LC_11_15_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance6.periodCounter_13_LC_11_15_5  (
            .in0(N__21421),
            .in1(N__23030),
            .in2(_gnd_net_),
            .in3(N__20412),
            .lcout(\PWMInstance6.periodCounterZ0Z_13 ),
            .ltout(),
            .carryin(\PWMInstance6.un1_periodCounter_2_cry_12 ),
            .carryout(\PWMInstance6.un1_periodCounter_2_cry_13 ),
            .clk(N__38562),
            .ce(),
            .sr(N__35296));
    defparam \PWMInstance6.periodCounter_14_LC_11_15_6 .C_ON=1'b1;
    defparam \PWMInstance6.periodCounter_14_LC_11_15_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.periodCounter_14_LC_11_15_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance6.periodCounter_14_LC_11_15_6  (
            .in0(_gnd_net_),
            .in1(N__23175),
            .in2(_gnd_net_),
            .in3(N__20409),
            .lcout(\PWMInstance6.periodCounterZ0Z_14 ),
            .ltout(),
            .carryin(\PWMInstance6.un1_periodCounter_2_cry_13 ),
            .carryout(\PWMInstance6.un1_periodCounter_2_cry_14 ),
            .clk(N__38562),
            .ce(),
            .sr(N__35296));
    defparam \PWMInstance6.periodCounter_15_LC_11_15_7 .C_ON=1'b1;
    defparam \PWMInstance6.periodCounter_15_LC_11_15_7 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.periodCounter_15_LC_11_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance6.periodCounter_15_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(N__23196),
            .in2(_gnd_net_),
            .in3(N__20406),
            .lcout(\PWMInstance6.periodCounterZ0Z_15 ),
            .ltout(),
            .carryin(\PWMInstance6.un1_periodCounter_2_cry_14 ),
            .carryout(\PWMInstance6.un1_periodCounter_2_cry_15 ),
            .clk(N__38562),
            .ce(),
            .sr(N__35296));
    defparam \PWMInstance6.periodCounter_16_LC_11_16_0 .C_ON=1'b0;
    defparam \PWMInstance6.periodCounter_16_LC_11_16_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.periodCounter_16_LC_11_16_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance6.periodCounter_16_LC_11_16_0  (
            .in0(N__21413),
            .in1(N__20923),
            .in2(_gnd_net_),
            .in3(N__20403),
            .lcout(\PWMInstance6.periodCounterZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38555),
            .ce(),
            .sr(N__35294));
    defparam \QuadInstance3.delayedCh_A_0_LC_12_1_3 .C_ON=1'b0;
    defparam \QuadInstance3.delayedCh_A_0_LC_12_1_3 .SEQ_MODE=4'b1000;
    defparam \QuadInstance3.delayedCh_A_0_LC_12_1_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance3.delayedCh_A_0_LC_12_1_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20400),
            .lcout(\QuadInstance3.delayedCh_AZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38702),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_RNIKINB1_14_LC_12_2_1 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_RNIKINB1_14_LC_12_2_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNIKINB1_14_LC_12_2_1 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \QuadInstance6.Quad_RNIKINB1_14_LC_12_2_1  (
            .in0(N__22791),
            .in1(N__22634),
            .in2(N__20562),
            .in3(N__22562),
            .lcout(\QuadInstance6.Quad_RNIKINB1Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_RNO_0_15_LC_12_3_6 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_RNO_0_15_LC_12_3_6 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNO_0_15_LC_12_3_6 .LUT_INIT=16'b0100101111110000;
    LogicCell40 \QuadInstance6.Quad_RNO_0_15_LC_12_3_6  (
            .in0(N__22792),
            .in1(N__22635),
            .in2(N__24273),
            .in3(N__22563),
            .lcout(\QuadInstance6.un1_Quad_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_5_LC_12_4_0 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_5_LC_12_4_0 .SEQ_MODE=4'b1000;
    defparam \QuadInstance1.Quad_5_LC_12_4_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \QuadInstance1.Quad_5_LC_12_4_0  (
            .in0(N__24100),
            .in1(N__21591),
            .in2(_gnd_net_),
            .in3(N__36371),
            .lcout(dataRead1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38680),
            .ce(),
            .sr(N__35693));
    defparam \QuadInstance2.Quad_5_LC_12_4_1 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_5_LC_12_4_1 .SEQ_MODE=4'b1000;
    defparam \QuadInstance2.Quad_5_LC_12_4_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \QuadInstance2.Quad_5_LC_12_4_1  (
            .in0(N__22191),
            .in1(_gnd_net_),
            .in2(N__36378),
            .in3(N__20370),
            .lcout(dataRead2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38680),
            .ce(),
            .sr(N__35693));
    defparam \QuadInstance6.Quad_7_LC_12_4_2 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_7_LC_12_4_2 .SEQ_MODE=4'b1000;
    defparam \QuadInstance6.Quad_7_LC_12_4_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \QuadInstance6.Quad_7_LC_12_4_2  (
            .in0(N__22794),
            .in1(_gnd_net_),
            .in2(N__29443),
            .in3(N__20499),
            .lcout(dataRead6_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38680),
            .ce(),
            .sr(N__35693));
    defparam \QuadInstance5.Quad_5_LC_12_4_3 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_5_LC_12_4_3 .SEQ_MODE=4'b1000;
    defparam \QuadInstance5.Quad_5_LC_12_4_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance5.Quad_5_LC_12_4_3  (
            .in0(N__36369),
            .in1(N__25795),
            .in2(_gnd_net_),
            .in3(N__20457),
            .lcout(dataRead5_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38680),
            .ce(),
            .sr(N__35693));
    defparam \QuadInstance6.Quad_5_LC_12_4_4 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_5_LC_12_4_4 .SEQ_MODE=4'b1000;
    defparam \QuadInstance6.Quad_5_LC_12_4_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance6.Quad_5_LC_12_4_4  (
            .in0(N__22793),
            .in1(N__36372),
            .in2(_gnd_net_),
            .in3(N__20517),
            .lcout(dataRead6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38680),
            .ce(),
            .sr(N__35693));
    defparam \QuadInstance7.Quad_5_LC_12_4_5 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_5_LC_12_4_5 .SEQ_MODE=4'b1000;
    defparam \QuadInstance7.Quad_5_LC_12_4_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance7.Quad_5_LC_12_4_5  (
            .in0(N__36370),
            .in1(N__26053),
            .in2(_gnd_net_),
            .in3(N__20445),
            .lcout(dataRead7_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38680),
            .ce(),
            .sr(N__35693));
    defparam \QuadInstance1.Quad_6_LC_12_4_6 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_6_LC_12_4_6 .SEQ_MODE=4'b1000;
    defparam \QuadInstance1.Quad_6_LC_12_4_6 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \QuadInstance1.Quad_6_LC_12_4_6  (
            .in0(N__24101),
            .in1(N__31111),
            .in2(N__21579),
            .in3(_gnd_net_),
            .lcout(dataRead1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38680),
            .ce(),
            .sr(N__35693));
    defparam \QuadInstance6.Quad_3_LC_12_4_7 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_3_LC_12_4_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance6.Quad_3_LC_12_4_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance6.Quad_3_LC_12_4_7  (
            .in0(N__32083),
            .in1(N__22795),
            .in2(_gnd_net_),
            .in3(N__20421),
            .lcout(dataRead6_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38680),
            .ce(),
            .sr(N__35693));
    defparam \QuadInstance6.un1_Quad_cry_0_c_LC_12_5_0 .C_ON=1'b1;
    defparam \QuadInstance6.un1_Quad_cry_0_c_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.un1_Quad_cry_0_c_LC_12_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \QuadInstance6.un1_Quad_cry_0_c_LC_12_5_0  (
            .in0(_gnd_net_),
            .in1(N__22555),
            .in2(N__30810),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_5_0_),
            .carryout(\QuadInstance6.un1_Quad_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_RNO_0_1_LC_12_5_1 .C_ON=1'b1;
    defparam \QuadInstance6.Quad_RNO_0_1_LC_12_5_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNO_0_1_LC_12_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance6.Quad_RNO_0_1_LC_12_5_1  (
            .in0(_gnd_net_),
            .in1(N__23783),
            .in2(N__20703),
            .in3(N__20433),
            .lcout(\QuadInstance6.Quad_RNO_0_5_1 ),
            .ltout(),
            .carryin(\QuadInstance6.un1_Quad_cry_0 ),
            .carryout(\QuadInstance6.un1_Quad_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_RNO_0_2_LC_12_5_2 .C_ON=1'b1;
    defparam \QuadInstance6.Quad_RNO_0_2_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNO_0_2_LC_12_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance6.Quad_RNO_0_2_LC_12_5_2  (
            .in0(_gnd_net_),
            .in1(N__30346),
            .in2(N__20688),
            .in3(N__20424),
            .lcout(\QuadInstance6.Quad_RNO_0_6_2 ),
            .ltout(),
            .carryin(\QuadInstance6.un1_Quad_cry_1 ),
            .carryout(\QuadInstance6.un1_Quad_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_RNO_0_3_LC_12_5_3 .C_ON=1'b1;
    defparam \QuadInstance6.Quad_RNO_0_3_LC_12_5_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNO_0_3_LC_12_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance6.Quad_RNO_0_3_LC_12_5_3  (
            .in0(_gnd_net_),
            .in1(N__27796),
            .in2(N__20664),
            .in3(N__20415),
            .lcout(\QuadInstance6.Quad_RNO_0_6_3 ),
            .ltout(),
            .carryin(\QuadInstance6.un1_Quad_cry_2 ),
            .carryout(\QuadInstance6.un1_Quad_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_RNO_0_4_LC_12_5_4 .C_ON=1'b1;
    defparam \QuadInstance6.Quad_RNO_0_4_LC_12_5_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNO_0_4_LC_12_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance6.Quad_RNO_0_4_LC_12_5_4  (
            .in0(_gnd_net_),
            .in1(N__21500),
            .in2(N__20784),
            .in3(N__20520),
            .lcout(\QuadInstance6.Quad_RNO_0_6_4 ),
            .ltout(),
            .carryin(\QuadInstance6.un1_Quad_cry_3 ),
            .carryout(\QuadInstance6.un1_Quad_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_RNO_0_5_LC_12_5_5 .C_ON=1'b1;
    defparam \QuadInstance6.Quad_RNO_0_5_LC_12_5_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNO_0_5_LC_12_5_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance6.Quad_RNO_0_5_LC_12_5_5  (
            .in0(_gnd_net_),
            .in1(N__36766),
            .in2(N__20652),
            .in3(N__20511),
            .lcout(\QuadInstance6.Quad_RNO_0_6_5 ),
            .ltout(),
            .carryin(\QuadInstance6.un1_Quad_cry_4 ),
            .carryout(\QuadInstance6.un1_Quad_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_RNO_0_6_LC_12_5_6 .C_ON=1'b1;
    defparam \QuadInstance6.Quad_RNO_0_6_LC_12_5_6 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNO_0_6_LC_12_5_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance6.Quad_RNO_0_6_LC_12_5_6  (
            .in0(_gnd_net_),
            .in1(N__27724),
            .in2(N__20760),
            .in3(N__20502),
            .lcout(\QuadInstance6.Quad_RNO_0_6_6 ),
            .ltout(),
            .carryin(\QuadInstance6.un1_Quad_cry_5 ),
            .carryout(\QuadInstance6.un1_Quad_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_RNO_0_7_LC_12_5_7 .C_ON=1'b1;
    defparam \QuadInstance6.Quad_RNO_0_7_LC_12_5_7 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNO_0_7_LC_12_5_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance6.Quad_RNO_0_7_LC_12_5_7  (
            .in0(_gnd_net_),
            .in1(N__26287),
            .in2(N__20748),
            .in3(N__20493),
            .lcout(\QuadInstance6.Quad_RNO_0_6_7 ),
            .ltout(),
            .carryin(\QuadInstance6.un1_Quad_cry_6 ),
            .carryout(\QuadInstance6.un1_Quad_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_RNO_0_8_LC_12_6_0 .C_ON=1'b1;
    defparam \QuadInstance6.Quad_RNO_0_8_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNO_0_8_LC_12_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance6.Quad_RNO_0_8_LC_12_6_0  (
            .in0(_gnd_net_),
            .in1(N__37783),
            .in2(N__20799),
            .in3(N__20484),
            .lcout(\QuadInstance6.Quad_RNO_0_6_8 ),
            .ltout(),
            .carryin(bfn_12_6_0_),
            .carryout(\QuadInstance6.un1_Quad_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_RNO_0_9_LC_12_6_1 .C_ON=1'b1;
    defparam \QuadInstance6.Quad_RNO_0_9_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNO_0_9_LC_12_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance6.Quad_RNO_0_9_LC_12_6_1  (
            .in0(_gnd_net_),
            .in1(N__25419),
            .in2(N__20640),
            .in3(N__20481),
            .lcout(\QuadInstance6.Quad_RNO_0_6_9 ),
            .ltout(),
            .carryin(\QuadInstance6.un1_Quad_cry_8 ),
            .carryout(\QuadInstance6.un1_Quad_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_RNO_0_10_LC_12_6_2 .C_ON=1'b1;
    defparam \QuadInstance6.Quad_RNO_0_10_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNO_0_10_LC_12_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance6.Quad_RNO_0_10_LC_12_6_2  (
            .in0(_gnd_net_),
            .in1(N__34609),
            .in2(N__21702),
            .in3(N__20478),
            .lcout(\QuadInstance6.Quad_RNO_0_6_10 ),
            .ltout(),
            .carryin(\QuadInstance6.un1_Quad_cry_9 ),
            .carryout(\QuadInstance6.un1_Quad_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_RNO_0_11_LC_12_6_3 .C_ON=1'b1;
    defparam \QuadInstance6.Quad_RNO_0_11_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNO_0_11_LC_12_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance6.Quad_RNO_0_11_LC_12_6_3  (
            .in0(_gnd_net_),
            .in1(N__20830),
            .in2(N__20676),
            .in3(N__20469),
            .lcout(\QuadInstance6.Quad_RNO_0_6_11 ),
            .ltout(),
            .carryin(\QuadInstance6.un1_Quad_cry_10 ),
            .carryout(\QuadInstance6.un1_Quad_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_RNO_0_12_LC_12_6_4 .C_ON=1'b1;
    defparam \QuadInstance6.Quad_RNO_0_12_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNO_0_12_LC_12_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance6.Quad_RNO_0_12_LC_12_6_4  (
            .in0(_gnd_net_),
            .in1(N__22289),
            .in2(N__20772),
            .in3(N__20628),
            .lcout(\QuadInstance6.Quad_RNO_0_6_12 ),
            .ltout(),
            .carryin(\QuadInstance6.un1_Quad_cry_11 ),
            .carryout(\QuadInstance6.un1_Quad_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_RNO_0_13_LC_12_6_5 .C_ON=1'b1;
    defparam \QuadInstance6.Quad_RNO_0_13_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNO_0_13_LC_12_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance6.Quad_RNO_0_13_LC_12_6_5  (
            .in0(_gnd_net_),
            .in1(N__22476),
            .in2(N__22839),
            .in3(N__20616),
            .lcout(\QuadInstance6.Quad_RNO_0_6_13 ),
            .ltout(),
            .carryin(\QuadInstance6.un1_Quad_cry_12 ),
            .carryout(\QuadInstance6.un1_Quad_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_RNO_0_14_LC_12_6_6 .C_ON=1'b1;
    defparam \QuadInstance6.Quad_RNO_0_14_LC_12_6_6 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNO_0_14_LC_12_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance6.Quad_RNO_0_14_LC_12_6_6  (
            .in0(_gnd_net_),
            .in1(N__20613),
            .in2(N__20554),
            .in3(N__20604),
            .lcout(\QuadInstance6.Quad_RNO_0_6_14 ),
            .ltout(),
            .carryin(\QuadInstance6.un1_Quad_cry_13 ),
            .carryout(\QuadInstance6.un1_Quad_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_15_LC_12_6_7 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_15_LC_12_6_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance6.Quad_15_LC_12_6_7 .LUT_INIT=16'b1011000111100100;
    LogicCell40 \QuadInstance6.Quad_15_LC_12_6_7  (
            .in0(N__22783),
            .in1(N__20601),
            .in2(N__31895),
            .in3(N__20592),
            .lcout(dataRead6_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38663),
            .ce(),
            .sr(N__35706));
    defparam \QuadInstance1.Quad_10_LC_12_7_0 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_10_LC_12_7_0 .SEQ_MODE=4'b1000;
    defparam \QuadInstance1.Quad_10_LC_12_7_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance1.Quad_10_LC_12_7_0  (
            .in0(N__36133),
            .in1(N__24096),
            .in2(_gnd_net_),
            .in3(N__21684),
            .lcout(dataRead1_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38651),
            .ce(),
            .sr(N__35715));
    defparam \QuadInstance6.Quad_1_LC_12_7_1 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_1_LC_12_7_1 .SEQ_MODE=4'b1000;
    defparam \QuadInstance6.Quad_1_LC_12_7_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance6.Quad_1_LC_12_7_1  (
            .in0(N__22788),
            .in1(N__31247),
            .in2(_gnd_net_),
            .in3(N__20589),
            .lcout(dataRead6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38651),
            .ce(),
            .sr(N__35715));
    defparam \QuadInstance7.Quad_8_LC_12_7_2 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_8_LC_12_7_2 .SEQ_MODE=4'b1000;
    defparam \QuadInstance7.Quad_8_LC_12_7_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance7.Quad_8_LC_12_7_2  (
            .in0(N__26054),
            .in1(N__28985),
            .in2(_gnd_net_),
            .in3(N__20580),
            .lcout(dataRead7_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38651),
            .ce(),
            .sr(N__35715));
    defparam \QuadInstance6.Quad_14_LC_12_7_3 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_14_LC_12_7_3 .SEQ_MODE=4'b1000;
    defparam \QuadInstance6.Quad_14_LC_12_7_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance6.Quad_14_LC_12_7_3  (
            .in0(N__22787),
            .in1(N__34374),
            .in2(_gnd_net_),
            .in3(N__20568),
            .lcout(dataRead6_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38651),
            .ce(),
            .sr(N__35715));
    defparam \QuadInstance6.Quad_10_LC_12_7_4 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_10_LC_12_7_4 .SEQ_MODE=4'b1000;
    defparam \QuadInstance6.Quad_10_LC_12_7_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance6.Quad_10_LC_12_7_4  (
            .in0(N__36134),
            .in1(N__22789),
            .in2(_gnd_net_),
            .in3(N__20526),
            .lcout(dataRead6_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38651),
            .ce(),
            .sr(N__35715));
    defparam \QuadInstance7.Quad_10_LC_12_7_5 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_10_LC_12_7_5 .SEQ_MODE=4'b1000;
    defparam \QuadInstance7.Quad_10_LC_12_7_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance7.Quad_10_LC_12_7_5  (
            .in0(N__36135),
            .in1(N__26055),
            .in2(_gnd_net_),
            .in3(N__20724),
            .lcout(dataRead7_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38651),
            .ce(),
            .sr(N__35715));
    defparam \QuadInstance1.Quad_14_LC_12_7_6 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_14_LC_12_7_6 .SEQ_MODE=4'b1000;
    defparam \QuadInstance1.Quad_14_LC_12_7_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance1.Quad_14_LC_12_7_6  (
            .in0(N__34373),
            .in1(N__24097),
            .in2(_gnd_net_),
            .in3(N__21657),
            .lcout(dataRead1_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38651),
            .ce(),
            .sr(N__35715));
    defparam \QuadInstance5.Quad_9_LC_12_7_7 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_9_LC_12_7_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance5.Quad_9_LC_12_7_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance5.Quad_9_LC_12_7_7  (
            .in0(N__28558),
            .in1(N__25802),
            .in2(_gnd_net_),
            .in3(N__20712),
            .lcout(dataRead5_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38651),
            .ce(),
            .sr(N__35715));
    defparam \QuadInstance6.Quad_RNI02A91_1_LC_12_8_0 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_RNI02A91_1_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNI02A91_1_LC_12_8_0 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance6.Quad_RNI02A91_1_LC_12_8_0  (
            .in0(N__23782),
            .in1(N__22704),
            .in2(N__22551),
            .in3(N__22604),
            .lcout(\QuadInstance6.Quad_RNI02A91Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.delayedCh_A_RNI4QLG_2_LC_12_8_1 .C_ON=1'b0;
    defparam \QuadInstance6.delayedCh_A_RNI4QLG_2_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.delayedCh_A_RNI4QLG_2_LC_12_8_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \QuadInstance6.delayedCh_A_RNI4QLG_2_LC_12_8_1  (
            .in0(N__22466),
            .in1(N__22862),
            .in2(N__21720),
            .in3(N__22845),
            .lcout(\QuadInstance6.count_enable ),
            .ltout(\QuadInstance6.count_enable_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_RNI13A91_2_LC_12_8_2 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_RNI13A91_2_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNI13A91_2_LC_12_8_2 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance6.Quad_RNI13A91_2_LC_12_8_2  (
            .in0(N__30354),
            .in1(N__22705),
            .in2(N__20691),
            .in3(N__22605),
            .lcout(\QuadInstance6.Quad_RNI13A91Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_RNIHFNB1_11_LC_12_8_3 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_RNIHFNB1_11_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNIHFNB1_11_LC_12_8_3 .LUT_INIT=16'b1100010011000100;
    LogicCell40 \QuadInstance6.Quad_RNIHFNB1_11_LC_12_8_3  (
            .in0(N__22610),
            .in1(N__22533),
            .in2(N__22758),
            .in3(N__20840),
            .lcout(\QuadInstance6.Quad_RNIHFNB1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_RNI24A91_3_LC_12_8_4 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_RNI24A91_3_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNI24A91_3_LC_12_8_4 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance6.Quad_RNI24A91_3_LC_12_8_4  (
            .in0(N__27812),
            .in1(N__22706),
            .in2(N__22552),
            .in3(N__22606),
            .lcout(\QuadInstance6.Quad_RNI24A91Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_RNI46A91_5_LC_12_8_5 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_RNI46A91_5_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNI46A91_5_LC_12_8_5 .LUT_INIT=16'b1111010100000000;
    LogicCell40 \QuadInstance6.Quad_RNI46A91_5_LC_12_8_5  (
            .in0(N__22607),
            .in1(N__36776),
            .in2(N__22756),
            .in3(N__22528),
            .lcout(\QuadInstance6.Quad_RNI46A91Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_RNI8AA91_9_LC_12_8_6 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_RNI8AA91_9_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNI8AA91_9_LC_12_8_6 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance6.Quad_RNI8AA91_9_LC_12_8_6  (
            .in0(N__25418),
            .in1(N__22710),
            .in2(N__22553),
            .in3(N__22609),
            .lcout(\QuadInstance6.Quad_RNI8AA91Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_RNI79A91_8_LC_12_8_7 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_RNI79A91_8_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNI79A91_8_LC_12_8_7 .LUT_INIT=16'b1111010100000000;
    LogicCell40 \QuadInstance6.Quad_RNI79A91_8_LC_12_8_7  (
            .in0(N__22608),
            .in1(N__37787),
            .in2(N__22757),
            .in3(N__22529),
            .lcout(\QuadInstance6.Quad_RNI79A91Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.delayedCh_B_RNI0PFF_2_LC_12_9_0 .C_ON=1'b0;
    defparam \QuadInstance6.delayedCh_B_RNI0PFF_2_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.delayedCh_B_RNI0PFF_2_LC_12_9_0 .LUT_INIT=16'b0000110011000000;
    LogicCell40 \QuadInstance6.delayedCh_B_RNI0PFF_2_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(N__34469),
            .in2(N__21719),
            .in3(N__22861),
            .lcout(\QuadInstance6.un1_count_enable_i_a2_0_1 ),
            .ltout(\QuadInstance6.un1_count_enable_i_a2_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_RNI35A91_4_LC_12_9_1 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_RNI35A91_4_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNI35A91_4_LC_12_9_1 .LUT_INIT=16'b1100111100000000;
    LogicCell40 \QuadInstance6.Quad_RNI35A91_4_LC_12_9_1  (
            .in0(N__21504),
            .in1(N__22717),
            .in2(N__20787),
            .in3(N__22534),
            .lcout(\QuadInstance6.Quad_RNI35A91Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.delayedCh_A_1_LC_12_9_2 .C_ON=1'b0;
    defparam \QuadInstance6.delayedCh_A_1_LC_12_9_2 .SEQ_MODE=4'b1000;
    defparam \QuadInstance6.delayedCh_A_1_LC_12_9_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \QuadInstance6.delayedCh_A_1_LC_12_9_2  (
            .in0(N__21111),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\QuadInstance6.delayedCh_AZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38632),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_RNIIGNB1_12_LC_12_9_3 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_RNIIGNB1_12_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNIIGNB1_12_LC_12_9_3 .LUT_INIT=16'b1100111100000000;
    LogicCell40 \QuadInstance6.Quad_RNIIGNB1_12_LC_12_9_3  (
            .in0(N__22282),
            .in1(N__22720),
            .in2(N__22631),
            .in3(N__22539),
            .lcout(\QuadInstance6.Quad_RNIIGNB1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_RNI57A91_6_LC_12_9_4 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_RNI57A91_6_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNI57A91_6_LC_12_9_4 .LUT_INIT=16'b1010000011110000;
    LogicCell40 \QuadInstance6.Quad_RNI57A91_6_LC_12_9_4  (
            .in0(N__22719),
            .in1(N__27740),
            .in2(N__22554),
            .in3(N__22614),
            .lcout(\QuadInstance6.Quad_RNI57A91Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_RNI68A91_7_LC_12_9_5 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_RNI68A91_7_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNI68A91_7_LC_12_9_5 .LUT_INIT=16'b1100111100000000;
    LogicCell40 \QuadInstance6.Quad_RNI68A91_7_LC_12_9_5  (
            .in0(N__26303),
            .in1(N__22718),
            .in2(N__22630),
            .in3(N__22538),
            .lcout(\QuadInstance6.Quad_RNI68A91Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_1_13_LC_12_9_6.C_ON=1'b0;
    defparam OutReg_ess_RNO_1_13_LC_12_9_6.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_1_13_LC_12_9_6.LUT_INIT=16'b1101100001010101;
    LogicCell40 OutReg_ess_RNO_1_13_LC_12_9_6 (
            .in0(N__20736),
            .in1(N__22822),
            .in2(N__26107),
            .in3(N__37748),
            .lcout(OutReg_ess_RNO_1Z0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam quadWrite_6_LC_12_9_7.C_ON=1'b0;
    defparam quadWrite_6_LC_12_9_7.SEQ_MODE=4'b1000;
    defparam quadWrite_6_LC_12_9_7.LUT_INIT=16'b1000000000000000;
    LogicCell40 quadWrite_6_LC_12_9_7 (
            .in0(N__33826),
            .in1(N__33599),
            .in2(N__33467),
            .in3(N__33203),
            .lcout(quadWriteZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38632),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_1_11_LC_12_10_0.C_ON=1'b0;
    defparam OutReg_ess_RNO_1_11_LC_12_10_0.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_1_11_LC_12_10_0.LUT_INIT=16'b1110010001010101;
    LogicCell40 OutReg_ess_RNO_1_11_LC_12_10_0 (
            .in0(N__22395),
            .in1(N__20876),
            .in2(N__20844),
            .in3(N__32839),
            .lcout(),
            .ltout(OutReg_ess_RNO_1Z0Z_11_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_0_11_LC_12_10_1.C_ON=1'b0;
    defparam OutReg_ess_RNO_0_11_LC_12_10_1.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_0_11_LC_12_10_1.LUT_INIT=16'b1111001111000000;
    LogicCell40 OutReg_ess_RNO_0_11_LC_12_10_1 (
            .in0(_gnd_net_),
            .in1(N__37560),
            .in2(N__20817),
            .in3(N__20814),
            .lcout(),
            .ltout(OutReg_ess_RNO_0Z0Z_11_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_11_LC_12_10_2.C_ON=1'b0;
    defparam OutReg_ess_11_LC_12_10_2.SEQ_MODE=4'b1001;
    defparam OutReg_ess_11_LC_12_10_2.LUT_INIT=16'b1010101010111000;
    LogicCell40 OutReg_ess_11_LC_12_10_2 (
            .in0(N__34911),
            .in1(N__38883),
            .in2(N__20808),
            .in3(N__37394),
            .lcout(OutRegZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38619),
            .ce(N__37251),
            .sr(N__37133));
    defparam OutReg_ess_13_LC_12_10_5.C_ON=1'b0;
    defparam OutReg_ess_13_LC_12_10_5.SEQ_MODE=4'b1001;
    defparam OutReg_ess_13_LC_12_10_5.LUT_INIT=16'b1111111000000100;
    LogicCell40 OutReg_ess_13_LC_12_10_5 (
            .in0(N__37395),
            .in1(N__20805),
            .in2(N__38911),
            .in3(N__22929),
            .lcout(OutRegZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38619),
            .ce(N__37251),
            .sr(N__37133));
    defparam dataWrite_0_LC_12_11_0.C_ON=1'b0;
    defparam dataWrite_0_LC_12_11_0.SEQ_MODE=4'b1000;
    defparam dataWrite_0_LC_12_11_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 dataWrite_0_LC_12_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38157),
            .lcout(dataWriteZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38610),
            .ce(N__24461),
            .sr(_gnd_net_));
    defparam dataWrite_1_LC_12_11_1.C_ON=1'b0;
    defparam dataWrite_1_LC_12_11_1.SEQ_MODE=4'b1000;
    defparam dataWrite_1_LC_12_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 dataWrite_1_LC_12_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37563),
            .lcout(dataWriteZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38610),
            .ce(N__24461),
            .sr(_gnd_net_));
    defparam dataWrite_10_LC_12_11_2.C_ON=1'b0;
    defparam dataWrite_10_LC_12_11_2.SEQ_MODE=4'b1000;
    defparam dataWrite_10_LC_12_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 dataWrite_10_LC_12_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22887),
            .lcout(dataWriteZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38610),
            .ce(N__24461),
            .sr(_gnd_net_));
    defparam dataWrite_11_LC_12_11_3.C_ON=1'b0;
    defparam dataWrite_11_LC_12_11_3.SEQ_MODE=4'b1000;
    defparam dataWrite_11_LC_12_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 dataWrite_11_LC_12_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22875),
            .lcout(dataWriteZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38610),
            .ce(N__24461),
            .sr(_gnd_net_));
    defparam dataWrite_12_LC_12_11_4.C_ON=1'b0;
    defparam dataWrite_12_LC_12_11_4.SEQ_MODE=4'b1000;
    defparam dataWrite_12_LC_12_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 dataWrite_12_LC_12_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22923),
            .lcout(dataWriteZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38610),
            .ce(N__24461),
            .sr(_gnd_net_));
    defparam dataWrite_13_LC_12_11_5.C_ON=1'b0;
    defparam dataWrite_13_LC_12_11_5.SEQ_MODE=4'b1000;
    defparam dataWrite_13_LC_12_11_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 dataWrite_13_LC_12_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22911),
            .lcout(dataWriteZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38610),
            .ce(N__24461),
            .sr(_gnd_net_));
    defparam dataWrite_14_LC_12_11_6.C_ON=1'b0;
    defparam dataWrite_14_LC_12_11_6.SEQ_MODE=4'b1000;
    defparam dataWrite_14_LC_12_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 dataWrite_14_LC_12_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22898),
            .lcout(dataWriteZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38610),
            .ce(N__24461),
            .sr(_gnd_net_));
    defparam dataWrite_15_LC_12_11_7.C_ON=1'b0;
    defparam dataWrite_15_LC_12_11_7.SEQ_MODE=4'b1000;
    defparam dataWrite_15_LC_12_11_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 dataWrite_15_LC_12_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20889),
            .lcout(dataWriteZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38610),
            .ce(N__24461),
            .sr(_gnd_net_));
    defparam data_received_esr_18_LC_12_12_0.C_ON=1'b0;
    defparam data_received_esr_18_LC_12_12_0.SEQ_MODE=4'b1000;
    defparam data_received_esr_18_LC_12_12_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 data_received_esr_18_LC_12_12_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20901),
            .lcout(data_receivedZ0Z_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38598),
            .ce(N__26181),
            .sr(N__26151));
    defparam data_received_esr_19_LC_12_12_1.C_ON=1'b0;
    defparam data_received_esr_19_LC_12_12_1.SEQ_MODE=4'b1000;
    defparam data_received_esr_19_LC_12_12_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 data_received_esr_19_LC_12_12_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20907),
            .lcout(data_receivedZ0Z_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38598),
            .ce(N__26181),
            .sr(N__26151));
    defparam data_received_esr_20_LC_12_12_2.C_ON=1'b0;
    defparam data_received_esr_20_LC_12_12_2.SEQ_MODE=4'b1000;
    defparam data_received_esr_20_LC_12_12_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 data_received_esr_20_LC_12_12_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22995),
            .lcout(data_receivedZ0Z_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38598),
            .ce(N__26181),
            .sr(N__26151));
    defparam data_received_esr_17_LC_12_12_3.C_ON=1'b0;
    defparam data_received_esr_17_LC_12_12_3.SEQ_MODE=4'b1000;
    defparam data_received_esr_17_LC_12_12_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 data_received_esr_17_LC_12_12_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20895),
            .lcout(data_receivedZ0Z_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38598),
            .ce(N__26181),
            .sr(N__26151));
    defparam data_received_esr_16_LC_12_12_4.C_ON=1'b0;
    defparam data_received_esr_16_LC_12_12_4.SEQ_MODE=4'b1000;
    defparam data_received_esr_16_LC_12_12_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 data_received_esr_16_LC_12_12_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20888),
            .lcout(data_receivedZ0Z_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38598),
            .ce(N__26181),
            .sr(N__26151));
    defparam data_received_esr_15_LC_12_12_5.C_ON=1'b0;
    defparam data_received_esr_15_LC_12_12_5.SEQ_MODE=4'b1000;
    defparam data_received_esr_15_LC_12_12_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 data_received_esr_15_LC_12_12_5 (
            .in0(N__22899),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(data_receivedZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38598),
            .ce(N__26181),
            .sr(N__26151));
    defparam data_received_esr_3_LC_12_12_6.C_ON=1'b0;
    defparam data_received_esr_3_LC_12_12_6.SEQ_MODE=4'b1000;
    defparam data_received_esr_3_LC_12_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 data_received_esr_3_LC_12_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37764),
            .lcout(data_receivedZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38598),
            .ce(N__26181),
            .sr(N__26151));
    defparam data_received_esr_21_LC_12_12_7.C_ON=1'b0;
    defparam data_received_esr_21_LC_12_12_7.SEQ_MODE=4'b1000;
    defparam data_received_esr_21_LC_12_12_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 data_received_esr_21_LC_12_12_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33586),
            .lcout(data_receivedZ0Z_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38598),
            .ce(N__26181),
            .sr(N__26151));
    defparam \PWMInstance6.clkCount_0_LC_12_13_1 .C_ON=1'b0;
    defparam \PWMInstance6.clkCount_0_LC_12_13_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.clkCount_0_LC_12_13_1 .LUT_INIT=16'b1010101000010001;
    LogicCell40 \PWMInstance6.clkCount_0_LC_12_13_1  (
            .in0(N__20942),
            .in1(N__20969),
            .in2(_gnd_net_),
            .in3(N__20990),
            .lcout(\PWMInstance6.clkCountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38591),
            .ce(),
            .sr(N__35757));
    defparam \PWMInstance6.clkCount_1_LC_12_13_6 .C_ON=1'b0;
    defparam \PWMInstance6.clkCount_1_LC_12_13_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.clkCount_1_LC_12_13_6 .LUT_INIT=16'b1100001011000010;
    LogicCell40 \PWMInstance6.clkCount_1_LC_12_13_6  (
            .in0(N__20991),
            .in1(N__20943),
            .in2(N__20973),
            .in3(_gnd_net_),
            .lcout(\PWMInstance6.clkCountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38591),
            .ce(),
            .sr(N__35757));
    defparam \PWMInstance6.out_RNO_0_LC_12_14_0 .C_ON=1'b0;
    defparam \PWMInstance6.out_RNO_0_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance6.out_RNO_0_LC_12_14_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \PWMInstance6.out_RNO_0_LC_12_14_0  (
            .in0(N__20952),
            .in1(N__20989),
            .in2(N__20928),
            .in3(N__20968),
            .lcout(\PWMInstance6.un1_periodCounter12_1_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwmWrite_6_LC_12_14_1.C_ON=1'b0;
    defparam pwmWrite_6_LC_12_14_1.SEQ_MODE=4'b1000;
    defparam pwmWrite_6_LC_12_14_1.LUT_INIT=16'b0010000000000000;
    LogicCell40 pwmWrite_6_LC_12_14_1 (
            .in0(N__33192),
            .in1(N__33456),
            .in2(N__33637),
            .in3(N__33783),
            .lcout(pwmWriteZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38580),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance6.clkCount_RNIBCT4_0_LC_12_14_2 .C_ON=1'b0;
    defparam \PWMInstance6.clkCount_RNIBCT4_0_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \PWMInstance6.clkCount_RNIBCT4_0_LC_12_14_2 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \PWMInstance6.clkCount_RNIBCT4_0_LC_12_14_2  (
            .in0(N__20951),
            .in1(N__20988),
            .in2(_gnd_net_),
            .in3(N__20967),
            .lcout(\PWMInstance6.periodCounter12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwmWrite_fast_6_LC_12_14_3.C_ON=1'b0;
    defparam pwmWrite_fast_6_LC_12_14_3.SEQ_MODE=4'b1000;
    defparam pwmWrite_fast_6_LC_12_14_3.LUT_INIT=16'b0010000000000000;
    LogicCell40 pwmWrite_fast_6_LC_12_14_3 (
            .in0(N__33193),
            .in1(N__33457),
            .in2(N__33638),
            .in3(N__33784),
            .lcout(pwmWrite_fastZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38580),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance6.PWMPulseWidthCount_esr_ctle_15_LC_12_14_4 .C_ON=1'b0;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_ctle_15_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_ctle_15_LC_12_14_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \PWMInstance6.PWMPulseWidthCount_esr_ctle_15_LC_12_14_4  (
            .in0(N__35829),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20941),
            .lcout(\PWMInstance6.pwmWrite_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance6.periodCounter_RNIET9F_16_LC_12_14_5 .C_ON=1'b0;
    defparam \PWMInstance6.periodCounter_RNIET9F_16_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \PWMInstance6.periodCounter_RNIET9F_16_LC_12_14_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \PWMInstance6.periodCounter_RNIET9F_16_LC_12_14_5  (
            .in0(_gnd_net_),
            .in1(N__20924),
            .in2(_gnd_net_),
            .in3(N__21022),
            .lcout(),
            .ltout(\PWMInstance6.un1_periodCounter12_1_0_a2_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance6.periodCounter_RNI00H31_15_LC_12_14_6 .C_ON=1'b0;
    defparam \PWMInstance6.periodCounter_RNI00H31_15_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \PWMInstance6.periodCounter_RNI00H31_15_LC_12_14_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \PWMInstance6.periodCounter_RNI00H31_15_LC_12_14_6  (
            .in0(N__21073),
            .in1(N__23188),
            .in2(N__21165),
            .in3(N__21154),
            .lcout(\PWMInstance6.un1_periodCounter12_1_0_a2_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.delayedCh_A_0_LC_12_14_7 .C_ON=1'b0;
    defparam \QuadInstance6.delayedCh_A_0_LC_12_14_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance6.delayedCh_A_0_LC_12_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance6.delayedCh_A_0_LC_12_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21126),
            .lcout(\QuadInstance6.delayedCh_AZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38580),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance6.periodCounter_RNI23321_13_LC_12_15_0 .C_ON=1'b0;
    defparam \PWMInstance6.periodCounter_RNI23321_13_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance6.periodCounter_RNI23321_13_LC_12_15_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \PWMInstance6.periodCounter_RNI23321_13_LC_12_15_0  (
            .in0(N__21089),
            .in1(N__23026),
            .in2(N__21042),
            .in3(N__21245),
            .lcout(\PWMInstance6.un1_periodCounter12_1_0_a2_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_12_15_1 .C_ON=1'b0;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_12_15_1 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance6.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_12_15_1  (
            .in0(N__21048),
            .in1(N__21088),
            .in2(N__21075),
            .in3(N__21054),
            .lcout(\PWMInstance6.un1_PWMPulseWidthCount_0_I_1_c_RNO_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance6.PWMPulseWidthCount_esr_0_LC_12_15_2 .C_ON=1'b0;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_0_LC_12_15_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_0_LC_12_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance6.PWMPulseWidthCount_esr_0_LC_12_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31378),
            .lcout(\PWMInstance6.PWMPulseWidthCountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38570),
            .ce(N__24557),
            .sr(N__35769));
    defparam \PWMInstance6.PWMPulseWidthCount_esr_1_LC_12_15_3 .C_ON=1'b0;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_1_LC_12_15_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_1_LC_12_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance6.PWMPulseWidthCount_esr_1_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31257),
            .lcout(\PWMInstance6.PWMPulseWidthCountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38570),
            .ce(N__24557),
            .sr(N__35769));
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_12_15_4 .C_ON=1'b0;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_12_15_4 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \PWMInstance6.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_12_15_4  (
            .in0(N__21037),
            .in1(N__21006),
            .in2(N__21000),
            .in3(N__21023),
            .lcout(\PWMInstance6.un1_PWMPulseWidthCount_0_I_27_c_RNO_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance6.PWMPulseWidthCount_esr_6_LC_12_15_5 .C_ON=1'b0;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_6_LC_12_15_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_6_LC_12_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance6.PWMPulseWidthCount_esr_6_LC_12_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31119),
            .lcout(\PWMInstance6.PWMPulseWidthCountZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38570),
            .ce(N__24557),
            .sr(N__35769));
    defparam \PWMInstance6.PWMPulseWidthCount_esr_7_LC_12_15_6 .C_ON=1'b0;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_7_LC_12_15_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_7_LC_12_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance6.PWMPulseWidthCount_esr_7_LC_12_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29444),
            .lcout(\PWMInstance6.PWMPulseWidthCountZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38570),
            .ce(N__24557),
            .sr(N__35769));
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_12_15_7 .C_ON=1'b0;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_12_15_7 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \PWMInstance6.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_12_15_7  (
            .in0(N__22947),
            .in1(N__21244),
            .in2(N__21228),
            .in3(N__24570),
            .lcout(\PWMInstance6.un1_PWMPulseWidthCount_0_I_45_c_RNO_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_1_c_LC_12_16_0 .C_ON=1'b1;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_1_c_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_1_c_LC_12_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance6.un1_PWMPulseWidthCount_0_I_1_c_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(N__21207),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_16_0_),
            .carryout(\PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_9_c_LC_12_16_1 .C_ON=1'b1;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_9_c_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_9_c_LC_12_16_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance6.un1_PWMPulseWidthCount_0_I_9_c_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(N__32314),
            .in2(N__21201),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_0 ),
            .carryout(\PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_15_c_LC_12_16_2 .C_ON=1'b1;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_15_c_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_15_c_LC_12_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance6.un1_PWMPulseWidthCount_0_I_15_c_LC_12_16_2  (
            .in0(_gnd_net_),
            .in1(N__21189),
            .in2(N__32410),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_1 ),
            .carryout(\PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_27_c_LC_12_16_3 .C_ON=1'b1;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_27_c_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_27_c_LC_12_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance6.un1_PWMPulseWidthCount_0_I_27_c_LC_12_16_3  (
            .in0(_gnd_net_),
            .in1(N__32306),
            .in2(N__21180),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_2 ),
            .carryout(\PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_45_c_LC_12_16_4 .C_ON=1'b1;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_45_c_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_45_c_LC_12_16_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance6.un1_PWMPulseWidthCount_0_I_45_c_LC_12_16_4  (
            .in0(_gnd_net_),
            .in1(N__21171),
            .in2(N__32412),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_3 ),
            .carryout(\PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_33_c_LC_12_16_5 .C_ON=1'b1;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_33_c_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_33_c_LC_12_16_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance6.un1_PWMPulseWidthCount_0_I_33_c_LC_12_16_5  (
            .in0(_gnd_net_),
            .in1(N__32307),
            .in2(N__23076),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_4 ),
            .carryout(\PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_39_c_LC_12_16_6 .C_ON=1'b1;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_39_c_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_39_c_LC_12_16_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance6.un1_PWMPulseWidthCount_0_I_39_c_LC_12_16_6  (
            .in0(_gnd_net_),
            .in1(N__23004),
            .in2(N__32411),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_5 ),
            .carryout(\PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_21_c_LC_12_16_7 .C_ON=1'b1;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_21_c_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_21_c_LC_12_16_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance6.un1_PWMPulseWidthCount_0_I_21_c_LC_12_16_7  (
            .in0(_gnd_net_),
            .in1(N__32305),
            .in2(N__23154),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_6 ),
            .carryout(\PWMInstance6.un1_PWMPulseWidthCount_0_data_tmp_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance6.out_LC_12_17_0 .C_ON=1'b0;
    defparam \PWMInstance6.out_LC_12_17_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.out_LC_12_17_0 .LUT_INIT=16'b1111101011110010;
    LogicCell40 \PWMInstance6.out_LC_12_17_0  (
            .in0(N__21368),
            .in1(N__21435),
            .in2(N__21426),
            .in3(N__21381),
            .lcout(PWM6_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38556),
            .ce(),
            .sr(N__35781));
    defparam PWM5_obufLegalizeSB_DFF_LC_12_20_0.C_ON=1'b0;
    defparam PWM5_obufLegalizeSB_DFF_LC_12_20_0.SEQ_MODE=4'b1000;
    defparam PWM5_obufLegalizeSB_DFF_LC_12_20_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 PWM5_obufLegalizeSB_DFF_LC_12_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PWM5_obufLegalizeSB_DFFNet),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36932),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance2.delayedCh_A_0_LC_13_2_0 .C_ON=1'b0;
    defparam \QuadInstance2.delayedCh_A_0_LC_13_2_0 .SEQ_MODE=4'b1000;
    defparam \QuadInstance2.delayedCh_A_0_LC_13_2_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \QuadInstance2.delayedCh_A_0_LC_13_2_0  (
            .in0(N__21351),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\QuadInstance2.delayedCh_AZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38703),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_1_LC_13_3_6 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_1_LC_13_3_6 .SEQ_MODE=4'b1000;
    defparam \QuadInstance1.Quad_1_LC_13_3_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance1.Quad_1_LC_13_3_6  (
            .in0(N__24059),
            .in1(N__31271),
            .in2(_gnd_net_),
            .in3(N__21645),
            .lcout(dataRead1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38695),
            .ce(),
            .sr(N__35694));
    defparam OutReg_ess_RNO_2_4_LC_13_4_0.C_ON=1'b0;
    defparam OutReg_ess_RNO_2_4_LC_13_4_0.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_2_4_LC_13_4_0.LUT_INIT=16'b1100000010111011;
    LogicCell40 OutReg_ess_RNO_2_4_LC_13_4_0 (
            .in0(N__21327),
            .in1(N__38153),
            .in2(N__23265),
            .in3(N__21252),
            .lcout(),
            .ltout(OutReg_ess_RNO_2Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_0_4_LC_13_4_1.C_ON=1'b0;
    defparam OutReg_ess_RNO_0_4_LC_13_4_1.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_0_4_LC_13_4_1.LUT_INIT=16'b1111110000110000;
    LogicCell40 OutReg_ess_RNO_0_4_LC_13_4_1 (
            .in0(_gnd_net_),
            .in1(N__37556),
            .in2(N__21300),
            .in3(N__21258),
            .lcout(OutReg_ess_RNO_0Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_3_4_LC_13_4_2.C_ON=1'b0;
    defparam OutReg_ess_RNO_3_4_LC_13_4_2.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_3_4_LC_13_4_2.LUT_INIT=16'b0101001001010111;
    LogicCell40 OutReg_ess_RNO_3_4_LC_13_4_2 (
            .in0(N__34763),
            .in1(N__21838),
            .in2(N__34896),
            .in3(N__21295),
            .lcout(),
            .ltout(OutReg_0_4_i_m3_ns_1_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_1_4_LC_13_4_3.C_ON=1'b0;
    defparam OutReg_ess_RNO_1_4_LC_13_4_3.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_1_4_LC_13_4_3.LUT_INIT=16'b1010110000001111;
    LogicCell40 OutReg_ess_RNO_1_4_LC_13_4_3 (
            .in0(N__21496),
            .in1(N__21451),
            .in2(N__21261),
            .in3(N__37737),
            .lcout(OutReg_ess_RNO_1Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_4_4_LC_13_4_4.C_ON=1'b0;
    defparam OutReg_ess_RNO_4_4_LC_13_4_4.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_4_4_LC_13_4_4.LUT_INIT=16'b0011000100111101;
    LogicCell40 OutReg_ess_RNO_4_4_LC_13_4_4 (
            .in0(N__34153),
            .in1(N__28138),
            .in2(N__28017),
            .in3(N__27517),
            .lcout(OutReg_0_5_i_m3_ns_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.delayedCh_A_0_LC_13_4_6 .C_ON=1'b0;
    defparam \QuadInstance0.delayedCh_A_0_LC_13_4_6 .SEQ_MODE=4'b1000;
    defparam \QuadInstance0.delayedCh_A_0_LC_13_4_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance0.delayedCh_A_0_LC_13_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21540),
            .lcout(\QuadInstance0.delayedCh_AZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38689),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_4_LC_13_5_0 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_4_LC_13_5_0 .SEQ_MODE=4'b1000;
    defparam \QuadInstance0.Quad_4_LC_13_5_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance0.Quad_4_LC_13_5_0  (
            .in0(N__33128),
            .in1(N__36484),
            .in2(_gnd_net_),
            .in3(N__29847),
            .lcout(dataRead0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38681),
            .ce(),
            .sr(N__35707));
    defparam \QuadInstance1.Quad_4_LC_13_5_1 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_4_LC_13_5_1 .SEQ_MODE=4'b1000;
    defparam \QuadInstance1.Quad_4_LC_13_5_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance1.Quad_4_LC_13_5_1  (
            .in0(N__36485),
            .in1(N__24051),
            .in2(_gnd_net_),
            .in3(N__21600),
            .lcout(dataRead1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38681),
            .ce(),
            .sr(N__35707));
    defparam \QuadInstance4.Quad_1_LC_13_5_2 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_1_LC_13_5_2 .SEQ_MODE=4'b1000;
    defparam \QuadInstance4.Quad_1_LC_13_5_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance4.Quad_1_LC_13_5_2  (
            .in0(N__29658),
            .in1(N__31252),
            .in2(_gnd_net_),
            .in3(N__24951),
            .lcout(dataRead4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38681),
            .ce(),
            .sr(N__35707));
    defparam \QuadInstance4.Quad_4_LC_13_5_3 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_4_LC_13_5_3 .SEQ_MODE=4'b1000;
    defparam \QuadInstance4.Quad_4_LC_13_5_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance4.Quad_4_LC_13_5_3  (
            .in0(N__36486),
            .in1(N__29659),
            .in2(_gnd_net_),
            .in3(N__24930),
            .lcout(dataRead4_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38681),
            .ce(),
            .sr(N__35707));
    defparam \QuadInstance3.Quad_6_LC_13_5_4 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_6_LC_13_5_4 .SEQ_MODE=4'b1000;
    defparam \QuadInstance3.Quad_6_LC_13_5_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance3.Quad_6_LC_13_5_4  (
            .in0(N__31109),
            .in1(N__22020),
            .in2(_gnd_net_),
            .in3(N__21525),
            .lcout(dataRead3_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38681),
            .ce(),
            .sr(N__35707));
    defparam \QuadInstance6.Quad_4_LC_13_5_5 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_4_LC_13_5_5 .SEQ_MODE=4'b1000;
    defparam \QuadInstance6.Quad_4_LC_13_5_5 .LUT_INIT=16'b1011100010111000;
    LogicCell40 \QuadInstance6.Quad_4_LC_13_5_5  (
            .in0(N__36487),
            .in1(N__22806),
            .in2(N__21513),
            .in3(_gnd_net_),
            .lcout(dataRead6_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38681),
            .ce(),
            .sr(N__35707));
    defparam \QuadInstance7.Quad_4_LC_13_5_6 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_4_LC_13_5_6 .SEQ_MODE=4'b1000;
    defparam \QuadInstance7.Quad_4_LC_13_5_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance7.Quad_4_LC_13_5_6  (
            .in0(N__26043),
            .in1(N__36488),
            .in2(_gnd_net_),
            .in3(N__21477),
            .lcout(dataRead7_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38681),
            .ce(),
            .sr(N__35707));
    defparam \QuadInstance0.Quad_9_LC_13_5_7 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_9_LC_13_5_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance0.Quad_9_LC_13_5_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance0.Quad_9_LC_13_5_7  (
            .in0(N__28565),
            .in1(N__33129),
            .in2(_gnd_net_),
            .in3(N__30117),
            .lcout(dataRead0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38681),
            .ce(),
            .sr(N__35707));
    defparam \QuadInstance1.un1_Quad_cry_0_c_LC_13_6_0 .C_ON=1'b1;
    defparam \QuadInstance1.un1_Quad_cry_0_c_LC_13_6_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.un1_Quad_cry_0_c_LC_13_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \QuadInstance1.un1_Quad_cry_0_c_LC_13_6_0  (
            .in0(_gnd_net_),
            .in1(N__24196),
            .in2(N__30943),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_6_0_),
            .carryout(\QuadInstance1.un1_Quad_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNO_0_1_LC_13_6_1 .C_ON=1'b1;
    defparam \QuadInstance1.Quad_RNO_0_1_LC_13_6_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNO_0_1_LC_13_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance1.Quad_RNO_0_1_LC_13_6_1  (
            .in0(_gnd_net_),
            .in1(N__23890),
            .in2(N__23538),
            .in3(N__21636),
            .lcout(\QuadInstance1.Quad_RNO_0_0_1 ),
            .ltout(),
            .carryin(\QuadInstance1.un1_Quad_cry_0 ),
            .carryout(\QuadInstance1.un1_Quad_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNO_0_2_LC_13_6_2 .C_ON=1'b1;
    defparam \QuadInstance1.Quad_RNO_0_2_LC_13_6_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNO_0_2_LC_13_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance1.Quad_RNO_0_2_LC_13_6_2  (
            .in0(_gnd_net_),
            .in1(N__30568),
            .in2(N__23676),
            .in3(N__21618),
            .lcout(\QuadInstance1.Quad_RNO_0_1_2 ),
            .ltout(),
            .carryin(\QuadInstance1.un1_Quad_cry_1 ),
            .carryout(\QuadInstance1.un1_Quad_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNO_0_3_LC_13_6_3 .C_ON=1'b1;
    defparam \QuadInstance1.Quad_RNO_0_3_LC_13_6_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNO_0_3_LC_13_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance1.Quad_RNO_0_3_LC_13_6_3  (
            .in0(_gnd_net_),
            .in1(N__27874),
            .in2(N__23667),
            .in3(N__21603),
            .lcout(\QuadInstance1.Quad_RNO_0_1_3 ),
            .ltout(),
            .carryin(\QuadInstance1.un1_Quad_cry_2 ),
            .carryout(\QuadInstance1.un1_Quad_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNO_0_4_LC_13_6_4 .C_ON=1'b1;
    defparam \QuadInstance1.Quad_RNO_0_4_LC_13_6_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNO_0_4_LC_13_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance1.Quad_RNO_0_4_LC_13_6_4  (
            .in0(_gnd_net_),
            .in1(N__23263),
            .in2(N__23241),
            .in3(N__21594),
            .lcout(\QuadInstance1.Quad_RNO_0_1_4 ),
            .ltout(),
            .carryin(\QuadInstance1.un1_Quad_cry_3 ),
            .carryout(\QuadInstance1.un1_Quad_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNO_0_5_LC_13_6_5 .C_ON=1'b1;
    defparam \QuadInstance1.Quad_RNO_0_5_LC_13_6_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNO_0_5_LC_13_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance1.Quad_RNO_0_5_LC_13_6_5  (
            .in0(_gnd_net_),
            .in1(N__36817),
            .in2(N__23520),
            .in3(N__21582),
            .lcout(\QuadInstance1.Quad_RNO_0_1_5 ),
            .ltout(),
            .carryin(\QuadInstance1.un1_Quad_cry_4 ),
            .carryout(\QuadInstance1.un1_Quad_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNO_0_6_LC_13_6_6 .C_ON=1'b1;
    defparam \QuadInstance1.Quad_RNO_0_6_LC_13_6_6 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNO_0_6_LC_13_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance1.Quad_RNO_0_6_LC_13_6_6  (
            .in0(_gnd_net_),
            .in1(N__25303),
            .in2(N__23529),
            .in3(N__21567),
            .lcout(\QuadInstance1.Quad_RNO_0_1_6 ),
            .ltout(),
            .carryin(\QuadInstance1.un1_Quad_cry_5 ),
            .carryout(\QuadInstance1.un1_Quad_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNO_0_7_LC_13_6_7 .C_ON=1'b1;
    defparam \QuadInstance1.Quad_RNO_0_7_LC_13_6_7 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNO_0_7_LC_13_6_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance1.Quad_RNO_0_7_LC_13_6_7  (
            .in0(_gnd_net_),
            .in1(N__25567),
            .in2(N__23685),
            .in3(N__21555),
            .lcout(\QuadInstance1.Quad_RNO_0_1_7 ),
            .ltout(),
            .carryin(\QuadInstance1.un1_Quad_cry_6 ),
            .carryout(\QuadInstance1.un1_Quad_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNO_0_8_LC_13_7_0 .C_ON=1'b1;
    defparam \QuadInstance1.Quad_RNO_0_8_LC_13_7_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNO_0_8_LC_13_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance1.Quad_RNO_0_8_LC_13_7_0  (
            .in0(_gnd_net_),
            .in1(N__37012),
            .in2(N__23634),
            .in3(N__21690),
            .lcout(\QuadInstance1.Quad_RNO_0_1_8 ),
            .ltout(),
            .carryin(bfn_13_7_0_),
            .carryout(\QuadInstance1.un1_Quad_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNO_0_9_LC_13_7_1 .C_ON=1'b1;
    defparam \QuadInstance1.Quad_RNO_0_9_LC_13_7_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNO_0_9_LC_13_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance1.Quad_RNO_0_9_LC_13_7_1  (
            .in0(_gnd_net_),
            .in1(N__25531),
            .in2(N__23481),
            .in3(N__21687),
            .lcout(\QuadInstance1.Quad_RNO_0_1_9 ),
            .ltout(),
            .carryin(\QuadInstance1.un1_Quad_cry_8 ),
            .carryout(\QuadInstance1.un1_Quad_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNO_0_10_LC_13_7_2 .C_ON=1'b1;
    defparam \QuadInstance1.Quad_RNO_0_10_LC_13_7_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNO_0_10_LC_13_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance1.Quad_RNO_0_10_LC_13_7_2  (
            .in0(_gnd_net_),
            .in1(N__35050),
            .in2(N__23472),
            .in3(N__21678),
            .lcout(\QuadInstance1.Quad_RNO_0_1_10 ),
            .ltout(),
            .carryin(\QuadInstance1.un1_Quad_cry_9 ),
            .carryout(\QuadInstance1.un1_Quad_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNO_0_11_LC_13_7_3 .C_ON=1'b1;
    defparam \QuadInstance1.Quad_RNO_0_11_LC_13_7_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNO_0_11_LC_13_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance1.Quad_RNO_0_11_LC_13_7_3  (
            .in0(_gnd_net_),
            .in1(N__23362),
            .in2(N__23340),
            .in3(N__21666),
            .lcout(\QuadInstance1.Quad_RNO_0_1_11 ),
            .ltout(),
            .carryin(\QuadInstance1.un1_Quad_cry_10 ),
            .carryout(\QuadInstance1.un1_Quad_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNO_0_12_LC_13_7_4 .C_ON=1'b1;
    defparam \QuadInstance1.Quad_RNO_0_12_LC_13_7_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNO_0_12_LC_13_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance1.Quad_RNO_0_12_LC_13_7_4  (
            .in0(_gnd_net_),
            .in1(N__24121),
            .in2(N__23658),
            .in3(N__21663),
            .lcout(\QuadInstance1.Quad_RNO_0_1_12 ),
            .ltout(),
            .carryin(\QuadInstance1.un1_Quad_cry_11 ),
            .carryout(\QuadInstance1.un1_Quad_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNO_0_13_LC_13_7_5 .C_ON=1'b1;
    defparam \QuadInstance1.Quad_RNO_0_13_LC_13_7_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNO_0_13_LC_13_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance1.Quad_RNO_0_13_LC_13_7_5  (
            .in0(_gnd_net_),
            .in1(N__23917),
            .in2(N__23649),
            .in3(N__21660),
            .lcout(\QuadInstance1.Quad_RNO_0_1_13 ),
            .ltout(),
            .carryin(\QuadInstance1.un1_Quad_cry_12 ),
            .carryout(\QuadInstance1.un1_Quad_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNO_0_14_LC_13_7_6 .C_ON=1'b1;
    defparam \QuadInstance1.Quad_RNO_0_14_LC_13_7_6 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNO_0_14_LC_13_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance1.Quad_RNO_0_14_LC_13_7_6  (
            .in0(_gnd_net_),
            .in1(N__23640),
            .in2(N__28189),
            .in3(N__21651),
            .lcout(\QuadInstance1.Quad_RNO_0_1_14 ),
            .ltout(),
            .carryin(\QuadInstance1.un1_Quad_cry_13 ),
            .carryout(\QuadInstance1.un1_Quad_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_15_LC_13_7_7 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_15_LC_13_7_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance1.Quad_15_LC_13_7_7 .LUT_INIT=16'b1101000111100010;
    LogicCell40 \QuadInstance1.Quad_15_LC_13_7_7  (
            .in0(N__23547),
            .in1(N__24050),
            .in2(N__31896),
            .in3(N__21648),
            .lcout(dataRead1_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38664),
            .ce(),
            .sr(N__35722));
    defparam \QuadInstance0.Quad_1_LC_13_8_0 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_1_LC_13_8_0 .SEQ_MODE=4'b1000;
    defparam \QuadInstance0.Quad_1_LC_13_8_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \QuadInstance0.Quad_1_LC_13_8_0  (
            .in0(N__31218),
            .in1(N__29892),
            .in2(_gnd_net_),
            .in3(N__33126),
            .lcout(dataRead0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38652),
            .ce(),
            .sr(N__35733));
    defparam \QuadInstance6.Quad_9_LC_13_8_1 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_9_LC_13_8_1 .SEQ_MODE=4'b1000;
    defparam \QuadInstance6.Quad_9_LC_13_8_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance6.Quad_9_LC_13_8_1  (
            .in0(N__22790),
            .in1(N__28528),
            .in2(_gnd_net_),
            .in3(N__22221),
            .lcout(dataRead6_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38652),
            .ce(),
            .sr(N__35733));
    defparam \QuadInstance2.Quad_1_LC_13_8_2 .C_ON=1'b0;
    defparam \QuadInstance2.Quad_1_LC_13_8_2 .SEQ_MODE=4'b1000;
    defparam \QuadInstance2.Quad_1_LC_13_8_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \QuadInstance2.Quad_1_LC_13_8_2  (
            .in0(N__31219),
            .in1(N__22209),
            .in2(_gnd_net_),
            .in3(N__22189),
            .lcout(dataRead2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38652),
            .ce(),
            .sr(N__35733));
    defparam \QuadInstance3.Quad_1_LC_13_8_3 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_1_LC_13_8_3 .SEQ_MODE=4'b1000;
    defparam \QuadInstance3.Quad_1_LC_13_8_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \QuadInstance3.Quad_1_LC_13_8_3  (
            .in0(N__22029),
            .in1(N__31220),
            .in2(_gnd_net_),
            .in3(N__22013),
            .lcout(dataRead3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38652),
            .ce(),
            .sr(N__35733));
    defparam \QuadInstance3.Quad_4_LC_13_8_4 .C_ON=1'b0;
    defparam \QuadInstance3.Quad_4_LC_13_8_4 .SEQ_MODE=4'b1000;
    defparam \QuadInstance3.Quad_4_LC_13_8_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \QuadInstance3.Quad_4_LC_13_8_4  (
            .in0(N__22012),
            .in1(_gnd_net_),
            .in2(N__36483),
            .in3(N__21855),
            .lcout(dataRead3_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38652),
            .ce(),
            .sr(N__35733));
    defparam \QuadInstance1.Quad_9_LC_13_8_5 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_9_LC_13_8_5 .SEQ_MODE=4'b1000;
    defparam \QuadInstance1.Quad_9_LC_13_8_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance1.Quad_9_LC_13_8_5  (
            .in0(N__24102),
            .in1(N__28527),
            .in2(_gnd_net_),
            .in3(N__21813),
            .lcout(dataRead1_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38652),
            .ce(),
            .sr(N__35733));
    defparam \QuadInstance6.Quad_0_LC_13_8_6 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_0_LC_13_8_6 .SEQ_MODE=4'b1000;
    defparam \QuadInstance6.Quad_0_LC_13_8_6 .LUT_INIT=16'b1011000111100100;
    LogicCell40 \QuadInstance6.Quad_0_LC_13_8_6  (
            .in0(N__22753),
            .in1(N__22550),
            .in2(N__31434),
            .in3(N__30799),
            .lcout(dataRead6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38652),
            .ce(),
            .sr(N__35733));
    defparam \QuadInstance7.Quad_0_LC_13_8_7 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_0_LC_13_8_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance7.Quad_0_LC_13_8_7 .LUT_INIT=16'b1100010111001010;
    LogicCell40 \QuadInstance7.Quad_0_LC_13_8_7  (
            .in0(N__30769),
            .in1(N__31407),
            .in2(N__26042),
            .in3(N__21807),
            .lcout(dataRead7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38652),
            .ce(),
            .sr(N__35733));
    defparam \QuadInstance6.delayedCh_B_2_LC_13_9_0 .C_ON=1'b0;
    defparam \QuadInstance6.delayedCh_B_2_LC_13_9_0 .SEQ_MODE=4'b1000;
    defparam \QuadInstance6.delayedCh_B_2_LC_13_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance6.delayedCh_B_2_LC_13_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22467),
            .lcout(\QuadInstance6.delayedCh_BZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38642),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_13_9_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_13_9_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_13_9_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_13_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_RNIGENB1_10_LC_13_9_2 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_RNIGENB1_10_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNIGENB1_10_LC_13_9_2 .LUT_INIT=16'b1100111100000000;
    LogicCell40 \QuadInstance6.Quad_RNIGENB1_10_LC_13_9_2  (
            .in0(N__34610),
            .in1(N__22721),
            .in2(N__22632),
            .in3(N__22548),
            .lcout(\QuadInstance6.Quad_RNIGENB1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.delayedCh_A_2_LC_13_9_3 .C_ON=1'b0;
    defparam \QuadInstance6.delayedCh_A_2_LC_13_9_3 .SEQ_MODE=4'b1000;
    defparam \QuadInstance6.delayedCh_A_2_LC_13_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance6.delayedCh_A_2_LC_13_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22863),
            .lcout(\QuadInstance6.delayedCh_AZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38642),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.Quad_RNIJHNB1_13_LC_13_9_4 .C_ON=1'b0;
    defparam \QuadInstance6.Quad_RNIJHNB1_13_LC_13_9_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance6.Quad_RNIJHNB1_13_LC_13_9_4 .LUT_INIT=16'b1100111100000000;
    LogicCell40 \QuadInstance6.Quad_RNIJHNB1_13_LC_13_9_4  (
            .in0(N__22838),
            .in1(N__22722),
            .in2(N__22633),
            .in3(N__22549),
            .lcout(\QuadInstance6.Quad_RNIJHNB1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.delayedCh_B_1_LC_13_9_6 .C_ON=1'b0;
    defparam \QuadInstance6.delayedCh_B_1_LC_13_9_6 .SEQ_MODE=4'b1000;
    defparam \QuadInstance6.delayedCh_B_1_LC_13_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance6.delayedCh_B_1_LC_13_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27108),
            .lcout(\QuadInstance6.delayedCh_BZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38642),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_3_11_LC_13_9_7.C_ON=1'b0;
    defparam OutReg_ess_RNO_3_11_LC_13_9_7.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_3_11_LC_13_9_7.LUT_INIT=16'b0000110100111101;
    LogicCell40 OutReg_ess_RNO_3_11_LC_13_9_7 (
            .in0(N__22450),
            .in1(N__34870),
            .in2(N__34772),
            .in3(N__22418),
            .lcout(OutReg_0_4_i_m3_i_m3_ns_1_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_esr_RNO_2_12_LC_13_10_0.C_ON=1'b0;
    defparam OutReg_esr_RNO_2_12_LC_13_10_0.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_2_12_LC_13_10_0.LUT_INIT=16'b1000100011110011;
    LogicCell40 OutReg_esr_RNO_2_12_LC_13_10_0 (
            .in0(N__24129),
            .in1(N__38138),
            .in2(N__22389),
            .in3(N__27624),
            .lcout(OutReg_esr_RNO_2Z0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_esr_RNO_3_12_LC_13_10_1.C_ON=1'b0;
    defparam OutReg_esr_RNO_3_12_LC_13_10_1.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_3_12_LC_13_10_1.LUT_INIT=16'b0000010110111011;
    LogicCell40 OutReg_esr_RNO_3_12_LC_13_10_1 (
            .in0(N__28126),
            .in1(N__22359),
            .in2(N__22331),
            .in3(N__28012),
            .lcout(),
            .ltout(OutReg_0_4_i_m3_ns_1_12_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_esr_RNO_1_12_LC_13_10_2.C_ON=1'b0;
    defparam OutReg_esr_RNO_1_12_LC_13_10_2.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_1_12_LC_13_10_2.LUT_INIT=16'b1010110000001111;
    LogicCell40 OutReg_esr_RNO_1_12_LC_13_10_2 (
            .in0(N__22293),
            .in1(N__22263),
            .in2(N__22233),
            .in3(N__37742),
            .lcout(),
            .ltout(OutReg_esr_RNO_1Z0Z_12_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_esr_RNO_0_12_LC_13_10_3.C_ON=1'b0;
    defparam OutReg_esr_RNO_0_12_LC_13_10_3.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_0_12_LC_13_10_3.LUT_INIT=16'b1111001111000000;
    LogicCell40 OutReg_esr_RNO_0_12_LC_13_10_3 (
            .in0(_gnd_net_),
            .in1(N__37559),
            .in2(N__22230),
            .in3(N__22227),
            .lcout(),
            .ltout(OutReg_esr_RNO_0Z0Z_12_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_esr_12_LC_13_10_4.C_ON=1'b0;
    defparam OutReg_esr_12_LC_13_10_4.SEQ_MODE=4'b1000;
    defparam OutReg_esr_12_LC_13_10_4.LUT_INIT=16'b1010101010111000;
    LogicCell40 OutReg_esr_12_LC_13_10_4 (
            .in0(N__22941),
            .in1(N__38951),
            .in2(N__22932),
            .in3(N__37388),
            .lcout(OutRegZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38633),
            .ce(N__37242),
            .sr(N__37130));
    defparam data_received_esr_13_LC_13_11_0.C_ON=1'b0;
    defparam data_received_esr_13_LC_13_11_0.SEQ_MODE=4'b1000;
    defparam data_received_esr_13_LC_13_11_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 data_received_esr_13_LC_13_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22922),
            .lcout(data_receivedZ0Z_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38620),
            .ce(N__26182),
            .sr(N__26152));
    defparam data_received_esr_10_LC_13_11_1.C_ON=1'b0;
    defparam data_received_esr_10_LC_13_11_1.SEQ_MODE=4'b1000;
    defparam data_received_esr_10_LC_13_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 data_received_esr_10_LC_13_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24474),
            .lcout(data_receivedZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38620),
            .ce(N__26182),
            .sr(N__26152));
    defparam data_received_esr_12_LC_13_11_2.C_ON=1'b0;
    defparam data_received_esr_12_LC_13_11_2.SEQ_MODE=4'b1000;
    defparam data_received_esr_12_LC_13_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 data_received_esr_12_LC_13_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22874),
            .lcout(data_receivedZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38620),
            .ce(N__26182),
            .sr(N__26152));
    defparam data_received_esr_14_LC_13_11_4.C_ON=1'b0;
    defparam data_received_esr_14_LC_13_11_4.SEQ_MODE=4'b1000;
    defparam data_received_esr_14_LC_13_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 data_received_esr_14_LC_13_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22910),
            .lcout(data_receivedZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38620),
            .ce(N__26182),
            .sr(N__26152));
    defparam data_received_esr_11_LC_13_11_6.C_ON=1'b0;
    defparam data_received_esr_11_LC_13_11_6.SEQ_MODE=4'b1000;
    defparam data_received_esr_11_LC_13_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 data_received_esr_11_LC_13_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22886),
            .lcout(data_receivedZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38620),
            .ce(N__26182),
            .sr(N__26152));
    defparam data_received_esr_23_LC_13_11_7.C_ON=1'b0;
    defparam data_received_esr_23_LC_13_11_7.SEQ_MODE=4'b1000;
    defparam data_received_esr_23_LC_13_11_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 data_received_esr_23_LC_13_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33283),
            .lcout(data_receivedZ0Z_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38620),
            .ce(N__26182),
            .sr(N__26152));
    defparam pwmWrite_3_LC_13_12_0.C_ON=1'b0;
    defparam pwmWrite_3_LC_13_12_0.SEQ_MODE=4'b1000;
    defparam pwmWrite_3_LC_13_12_0.LUT_INIT=16'b0000010000000000;
    LogicCell40 pwmWrite_3_LC_13_12_0 (
            .in0(N__33759),
            .in1(N__33557),
            .in2(N__33468),
            .in3(N__23391),
            .lcout(pwmWriteZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38611),
            .ce(),
            .sr(_gnd_net_));
    defparam data_received_esr_RNIMIH31_19_LC_13_12_1.C_ON=1'b0;
    defparam data_received_esr_RNIMIH31_19_LC_13_12_1.SEQ_MODE=4'b0000;
    defparam data_received_esr_RNIMIH31_19_LC_13_12_1.LUT_INIT=16'b0010000000000000;
    LogicCell40 data_received_esr_RNIMIH31_19_LC_13_12_1 (
            .in0(N__22994),
            .in1(N__37985),
            .in2(N__22980),
            .in3(N__39064),
            .lcout(data_received_esr_RNIMIH31Z0Z_19),
            .ltout(data_received_esr_RNIMIH31Z0Z_19_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwmWrite_fast_3_LC_13_12_2.C_ON=1'b0;
    defparam pwmWrite_fast_3_LC_13_12_2.SEQ_MODE=4'b1000;
    defparam pwmWrite_fast_3_LC_13_12_2.LUT_INIT=16'b0001000000000000;
    LogicCell40 pwmWrite_fast_3_LC_13_12_2 (
            .in0(N__33761),
            .in1(N__33459),
            .in2(N__22998),
            .in3(N__33559),
            .lcout(pwmWrite_fastZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38611),
            .ce(),
            .sr(_gnd_net_));
    defparam data_received_esr_RNIBPOR_23_LC_13_12_3.C_ON=1'b0;
    defparam data_received_esr_RNIBPOR_23_LC_13_12_3.SEQ_MODE=4'b0000;
    defparam data_received_esr_RNIBPOR_23_LC_13_12_3.LUT_INIT=16'b0010001000000000;
    LogicCell40 data_received_esr_RNIBPOR_23_LC_13_12_3 (
            .in0(N__22978),
            .in1(N__37986),
            .in2(_gnd_net_),
            .in3(N__39066),
            .lcout(N_870_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_received_esr_RNIMIH31_0_19_LC_13_12_5.C_ON=1'b0;
    defparam data_received_esr_RNIMIH31_0_19_LC_13_12_5.SEQ_MODE=4'b0000;
    defparam data_received_esr_RNIMIH31_0_19_LC_13_12_5.LUT_INIT=16'b0001000000000000;
    LogicCell40 data_received_esr_RNIMIH31_0_19_LC_13_12_5 (
            .in0(N__22993),
            .in1(N__37984),
            .in2(N__22979),
            .in3(N__39065),
            .lcout(data_received_esr_RNIMIH31_0Z0Z_19),
            .ltout(data_received_esr_RNIMIH31_0Z0Z_19_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwmWrite_fast_2_LC_13_12_6.C_ON=1'b0;
    defparam pwmWrite_fast_2_LC_13_12_6.SEQ_MODE=4'b1000;
    defparam pwmWrite_fast_2_LC_13_12_6.LUT_INIT=16'b0001000000000000;
    LogicCell40 pwmWrite_fast_2_LC_13_12_6 (
            .in0(N__33760),
            .in1(N__33458),
            .in2(N__22962),
            .in3(N__33558),
            .lcout(pwmWrite_fastZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38611),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance4.PWMPulseWidthCount_esr_0_LC_13_13_0 .C_ON=1'b0;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_0_LC_13_13_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_0_LC_13_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance4.PWMPulseWidthCount_esr_0_LC_13_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31382),
            .lcout(\PWMInstance4.PWMPulseWidthCountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38599),
            .ce(N__26958),
            .sr(N__35764));
    defparam \PWMInstance6.PWMPulseWidthCount_esr_13_LC_13_14_0 .C_ON=1'b0;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_13_LC_13_14_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_13_LC_13_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance6.PWMPulseWidthCount_esr_13_LC_13_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28677),
            .lcout(\PWMInstance6.PWMPulseWidthCountZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38592),
            .ce(N__24539),
            .sr(N__35770));
    defparam \PWMInstance6.PWMPulseWidthCount_esr_5_LC_13_14_1 .C_ON=1'b0;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_5_LC_13_14_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_5_LC_13_14_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \PWMInstance6.PWMPulseWidthCount_esr_5_LC_13_14_1  (
            .in0(_gnd_net_),
            .in1(N__36332),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PWMInstance6.PWMPulseWidthCountZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38592),
            .ce(N__24539),
            .sr(N__35770));
    defparam \PWMInstance6.PWMPulseWidthCount_esr_8_LC_13_14_2 .C_ON=1'b0;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_8_LC_13_14_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_8_LC_13_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance6.PWMPulseWidthCount_esr_8_LC_13_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28943),
            .lcout(\PWMInstance6.PWMPulseWidthCountZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38592),
            .ce(N__24539),
            .sr(N__35770));
    defparam \PWMInstance6.PWMPulseWidthCount_esr_11_LC_13_14_3 .C_ON=1'b0;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_11_LC_13_14_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_11_LC_13_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance6.PWMPulseWidthCount_esr_11_LC_13_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35994),
            .lcout(\PWMInstance6.PWMPulseWidthCountZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38592),
            .ce(N__24539),
            .sr(N__35770));
    defparam \PWMInstance6.PWMPulseWidthCount_esr_12_LC_13_14_6 .C_ON=1'b0;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_12_LC_13_14_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_12_LC_13_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance6.PWMPulseWidthCount_esr_12_LC_13_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28823),
            .lcout(\PWMInstance6.PWMPulseWidthCountZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38592),
            .ce(N__24539),
            .sr(N__35770));
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_13_15_0 .C_ON=1'b0;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_13_15_0 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance6.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_13_15_0  (
            .in0(N__23195),
            .in1(N__23145),
            .in2(N__23139),
            .in3(N__23174),
            .lcout(\PWMInstance6.un1_PWMPulseWidthCount_0_I_21_c_RNO_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance6.PWMPulseWidthCount_esr_14_LC_13_15_1 .C_ON=1'b0;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_14_LC_13_15_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_14_LC_13_15_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \PWMInstance6.PWMPulseWidthCount_esr_14_LC_13_15_1  (
            .in0(N__34394),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PWMInstance6.PWMPulseWidthCountZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38581),
            .ce(N__24558),
            .sr(N__35774));
    defparam \PWMInstance6.PWMPulseWidthCount_esr_15_LC_13_15_2 .C_ON=1'b0;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_15_LC_13_15_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_15_LC_13_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance6.PWMPulseWidthCount_esr_15_LC_13_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31857),
            .lcout(\PWMInstance6.PWMPulseWidthCountZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38581),
            .ce(N__24558),
            .sr(N__35774));
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_13_15_3 .C_ON=1'b0;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_13_15_3 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \PWMInstance6.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_13_15_3  (
            .in0(N__23130),
            .in1(N__23109),
            .in2(N__23103),
            .in3(N__23067),
            .lcout(\PWMInstance6.un1_PWMPulseWidthCount_0_I_33_c_RNO_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance6.PWMPulseWidthCount_esr_10_LC_13_15_4 .C_ON=1'b0;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_10_LC_13_15_4 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_10_LC_13_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance6.PWMPulseWidthCount_esr_10_LC_13_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36158),
            .lcout(\PWMInstance6.PWMPulseWidthCountZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38581),
            .ce(N__24558),
            .sr(N__35774));
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_13_15_6 .C_ON=1'b0;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_13_15_6 .SEQ_MODE=4'b0000;
    defparam \PWMInstance6.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_13_15_6 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance6.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_13_15_6  (
            .in0(N__23061),
            .in1(N__23055),
            .in2(N__23034),
            .in3(N__23010),
            .lcout(\PWMInstance6.un1_PWMPulseWidthCount_0_I_39_c_RNO_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance4.PWMPulseWidthCount_esr_12_LC_13_16_0 .C_ON=1'b0;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_12_LC_13_16_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_12_LC_13_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance4.PWMPulseWidthCount_esr_12_LC_13_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28854),
            .lcout(\PWMInstance4.PWMPulseWidthCountZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38571),
            .ce(N__26953),
            .sr(N__35782));
    defparam \PWMInstance4.PWMPulseWidthCount_esr_13_LC_13_16_1 .C_ON=1'b0;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_13_LC_13_16_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_13_LC_13_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance4.PWMPulseWidthCount_esr_13_LC_13_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28711),
            .lcout(\PWMInstance4.PWMPulseWidthCountZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38571),
            .ce(N__26953),
            .sr(N__35782));
    defparam \PWMInstance4.PWMPulseWidthCount_esr_8_LC_13_16_2 .C_ON=1'b0;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_8_LC_13_16_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_8_LC_13_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance4.PWMPulseWidthCount_esr_8_LC_13_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28976),
            .lcout(\PWMInstance4.PWMPulseWidthCountZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38571),
            .ce(N__26953),
            .sr(N__35782));
    defparam \PWMInstance4.PWMPulseWidthCount_esr_9_LC_13_16_3 .C_ON=1'b0;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_9_LC_13_16_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_9_LC_13_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance4.PWMPulseWidthCount_esr_9_LC_13_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28557),
            .lcout(\PWMInstance4.PWMPulseWidthCountZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38571),
            .ce(N__26953),
            .sr(N__35782));
    defparam \PWMInstance4.PWMPulseWidthCount_esr_3_LC_13_16_7 .C_ON=1'b0;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_3_LC_13_16_7 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_3_LC_13_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance4.PWMPulseWidthCount_esr_3_LC_13_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32043),
            .lcout(\PWMInstance4.PWMPulseWidthCountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38571),
            .ce(N__26953),
            .sr(N__35782));
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_13_17_0 .C_ON=1'b0;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_13_17_0 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance4.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_13_17_0  (
            .in0(N__23208),
            .in1(N__24652),
            .in2(N__24834),
            .in3(N__23214),
            .lcout(\PWMInstance4.un1_PWMPulseWidthCount_0_I_15_c_RNO_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance4.periodCounter_RNI3G5D_2_LC_13_17_1 .C_ON=1'b0;
    defparam \PWMInstance4.periodCounter_RNI3G5D_2_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance4.periodCounter_RNI3G5D_2_LC_13_17_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \PWMInstance4.periodCounter_RNI3G5D_2_LC_13_17_1  (
            .in0(_gnd_net_),
            .in1(N__24910),
            .in2(_gnd_net_),
            .in3(N__24694),
            .lcout(),
            .ltout(\PWMInstance4.un1_periodCounter12_1_0_a2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance4.periodCounter_RNIDRK61_4_LC_13_17_2 .C_ON=1'b0;
    defparam \PWMInstance4.periodCounter_RNIDRK61_4_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \PWMInstance4.periodCounter_RNIDRK61_4_LC_13_17_2 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \PWMInstance4.periodCounter_RNIDRK61_4_LC_13_17_2  (
            .in0(N__24745),
            .in1(N__24797),
            .in2(N__23217),
            .in3(N__24653),
            .lcout(\PWMInstance4.un1_periodCounter12_1_0_a2_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance4.PWMPulseWidthCount_esr_4_LC_13_17_3 .C_ON=1'b0;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_4_LC_13_17_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_4_LC_13_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance4.PWMPulseWidthCount_esr_4_LC_13_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36502),
            .lcout(\PWMInstance4.PWMPulseWidthCountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38563),
            .ce(N__26952),
            .sr(N__35786));
    defparam \PWMInstance4.PWMPulseWidthCount_esr_5_LC_13_17_4 .C_ON=1'b0;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_5_LC_13_17_4 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_5_LC_13_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance4.PWMPulseWidthCount_esr_5_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36362),
            .lcout(\PWMInstance4.PWMPulseWidthCountZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38563),
            .ce(N__26952),
            .sr(N__35786));
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_13_17_5 .C_ON=1'b0;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_13_17_5 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \PWMInstance4.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_13_17_5  (
            .in0(N__24796),
            .in1(N__23331),
            .in2(N__24776),
            .in3(N__23202),
            .lcout(\PWMInstance4.un1_PWMPulseWidthCount_0_I_33_c_RNO_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance4.PWMPulseWidthCount_esr_10_LC_13_17_6 .C_ON=1'b0;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_10_LC_13_17_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_10_LC_13_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance4.PWMPulseWidthCount_esr_10_LC_13_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36159),
            .lcout(\PWMInstance4.PWMPulseWidthCountZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38563),
            .ce(N__26952),
            .sr(N__35786));
    defparam \PWMInstance4.PWMPulseWidthCount_esr_11_LC_13_17_7 .C_ON=1'b0;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_11_LC_13_17_7 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_11_LC_13_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance4.PWMPulseWidthCount_esr_11_LC_13_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36014),
            .lcout(\PWMInstance4.PWMPulseWidthCountZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38563),
            .ce(N__26952),
            .sr(N__35786));
    defparam \QuadInstance2.delayedCh_B_0_LC_14_1_7 .C_ON=1'b0;
    defparam \QuadInstance2.delayedCh_B_0_LC_14_1_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance2.delayedCh_B_0_LC_14_1_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \QuadInstance2.delayedCh_B_0_LC_14_1_7  (
            .in0(N__23325),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\QuadInstance2.delayedCh_BZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38716),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.delayedCh_B_0_LC_14_2_7 .C_ON=1'b0;
    defparam \QuadInstance4.delayedCh_B_0_LC_14_2_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance4.delayedCh_B_0_LC_14_2_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \QuadInstance4.delayedCh_B_0_LC_14_2_7  (
            .in0(N__23295),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\QuadInstance4.delayedCh_BZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38710),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.delayedCh_A_0_LC_14_3_0 .C_ON=1'b0;
    defparam \QuadInstance4.delayedCh_A_0_LC_14_3_0 .SEQ_MODE=4'b1000;
    defparam \QuadInstance4.delayedCh_A_0_LC_14_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance4.delayedCh_A_0_LC_14_3_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23280),
            .lcout(\QuadInstance4.delayedCh_AZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38704),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.delayedCh_B_1_LC_14_3_5 .C_ON=1'b0;
    defparam \QuadInstance1.delayedCh_B_1_LC_14_3_5 .SEQ_MODE=4'b1000;
    defparam \QuadInstance1.delayedCh_B_1_LC_14_3_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance1.delayedCh_B_1_LC_14_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27072),
            .lcout(\QuadInstance1.delayedCh_BZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38704),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.delayedCh_B_2_LC_14_4_1 .C_ON=1'b0;
    defparam \QuadInstance1.delayedCh_B_2_LC_14_4_1 .SEQ_MODE=4'b1000;
    defparam \QuadInstance1.delayedCh_B_2_LC_14_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance1.delayedCh_B_2_LC_14_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23231),
            .lcout(\QuadInstance1.delayedCh_BZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38696),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.delayedCh_A_1_LC_14_4_6 .C_ON=1'b0;
    defparam \QuadInstance1.delayedCh_A_1_LC_14_4_6 .SEQ_MODE=4'b1000;
    defparam \QuadInstance1.delayedCh_A_1_LC_14_4_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance1.delayedCh_A_1_LC_14_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32118),
            .lcout(\QuadInstance1.delayedCh_AZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38696),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNIRK0O_4_LC_14_5_0 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_RNIRK0O_4_LC_14_5_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNIRK0O_4_LC_14_5_0 .LUT_INIT=16'b1111001100000000;
    LogicCell40 \QuadInstance1.Quad_RNIRK0O_4_LC_14_5_0  (
            .in0(N__23264),
            .in1(N__23580),
            .in2(N__24084),
            .in3(N__24180),
            .lcout(\QuadInstance1.Quad_RNIRK0OZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.delayedCh_A_RNIGDO2_2_LC_14_5_1 .C_ON=1'b0;
    defparam \QuadInstance1.delayedCh_A_RNIGDO2_2_LC_14_5_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.delayedCh_A_RNIGDO2_2_LC_14_5_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \QuadInstance1.delayedCh_A_RNIGDO2_2_LC_14_5_1  (
            .in0(N__23502),
            .in1(N__23492),
            .in2(N__23511),
            .in3(N__23232),
            .lcout(\QuadInstance1.count_enable ),
            .ltout(\QuadInstance1.count_enable_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNIOH0O_1_LC_14_5_2 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_RNIOH0O_1_LC_14_5_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNIOH0O_1_LC_14_5_2 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance1.Quad_RNIOH0O_1_LC_14_5_2  (
            .in0(N__23898),
            .in1(N__24004),
            .in2(N__23541),
            .in3(N__23579),
            .lcout(\QuadInstance1.Quad_RNIOH0OZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNITM0O_6_LC_14_5_3 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_RNITM0O_6_LC_14_5_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNITM0O_6_LC_14_5_3 .LUT_INIT=16'b1000101010001010;
    LogicCell40 \QuadInstance1.Quad_RNITM0O_6_LC_14_5_3  (
            .in0(N__24181),
            .in1(N__24052),
            .in2(N__23610),
            .in3(N__25311),
            .lcout(\QuadInstance1.Quad_RNITM0OZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNISL0O_5_LC_14_5_4 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_RNISL0O_5_LC_14_5_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNISL0O_5_LC_14_5_4 .LUT_INIT=16'b1111001100000000;
    LogicCell40 \QuadInstance1.Quad_RNISL0O_5_LC_14_5_4  (
            .in0(N__36827),
            .in1(N__23581),
            .in2(N__24085),
            .in3(N__24182),
            .lcout(\QuadInstance1.Quad_RNISL0OZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.delayedCh_A_2_LC_14_5_5 .C_ON=1'b0;
    defparam \QuadInstance1.delayedCh_A_2_LC_14_5_5 .SEQ_MODE=4'b1000;
    defparam \QuadInstance1.delayedCh_A_2_LC_14_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance1.delayedCh_A_2_LC_14_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23493),
            .lcout(\QuadInstance1.delayedCh_AZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38690),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.delayedCh_B_RNIM2H8_2_LC_14_5_7 .C_ON=1'b0;
    defparam \QuadInstance1.delayedCh_B_RNIM2H8_2_LC_14_5_7 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.delayedCh_B_RNIM2H8_2_LC_14_5_7 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \QuadInstance1.delayedCh_B_RNIM2H8_2_LC_14_5_7  (
            .in0(N__23501),
            .in1(N__34495),
            .in2(_gnd_net_),
            .in3(N__23491),
            .lcout(\QuadInstance1.un1_count_enable_i_a2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNI0Q0O_9_LC_14_6_0 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_RNI0Q0O_9_LC_14_6_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNI0Q0O_9_LC_14_6_0 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance1.Quad_RNI0Q0O_9_LC_14_6_0  (
            .in0(N__25545),
            .in1(N__24008),
            .in2(N__24198),
            .in3(N__23595),
            .lcout(\QuadInstance1.Quad_RNI0Q0OZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNI8P5D_10_LC_14_6_1 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_RNI8P5D_10_LC_14_6_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNI8P5D_10_LC_14_6_1 .LUT_INIT=16'b1010111100000000;
    LogicCell40 \QuadInstance1.Quad_RNI8P5D_10_LC_14_6_1  (
            .in0(N__24009),
            .in1(N__35061),
            .in2(N__23613),
            .in3(N__24178),
            .lcout(\QuadInstance1.Quad_RNI8P5DZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam quadWrite_1_LC_14_6_2.C_ON=1'b0;
    defparam quadWrite_1_LC_14_6_2.SEQ_MODE=4'b1000;
    defparam quadWrite_1_LC_14_6_2.LUT_INIT=16'b0001000000000000;
    LogicCell40 quadWrite_1_LC_14_6_2 (
            .in0(N__33858),
            .in1(N__33656),
            .in2(N__33448),
            .in3(N__23448),
            .lcout(quadWriteZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38682),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNI9Q5D_11_LC_14_6_3 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_RNI9Q5D_11_LC_14_6_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNI9Q5D_11_LC_14_6_3 .LUT_INIT=16'b1010111100000000;
    LogicCell40 \QuadInstance1.Quad_RNI9Q5D_11_LC_14_6_3  (
            .in0(N__24010),
            .in1(N__23370),
            .in2(N__23614),
            .in3(N__24179),
            .lcout(\QuadInstance1.Quad_RNI9Q5DZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_3_5_LC_14_6_4.C_ON=1'b0;
    defparam OutReg_ess_RNO_3_5_LC_14_6_4.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_3_5_LC_14_6_4.LUT_INIT=16'b0101001001010111;
    LogicCell40 OutReg_ess_RNO_3_5_LC_14_6_4 (
            .in0(N__34731),
            .in1(N__23734),
            .in2(N__34889),
            .in3(N__23710),
            .lcout(OutReg_0_4_i_m3_ns_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNIUN0O_7_LC_14_6_5 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_RNIUN0O_7_LC_14_6_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNIUN0O_7_LC_14_6_5 .LUT_INIT=16'b1010111100000000;
    LogicCell40 \QuadInstance1.Quad_RNIUN0O_7_LC_14_6_5  (
            .in0(N__24007),
            .in1(N__25568),
            .in2(N__23612),
            .in3(N__24174),
            .lcout(\QuadInstance1.Quad_RNIUN0OZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNIPI0O_2_LC_14_6_6 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_RNIPI0O_2_LC_14_6_6 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNIPI0O_2_LC_14_6_6 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance1.Quad_RNIPI0O_2_LC_14_6_6  (
            .in0(N__30569),
            .in1(N__24005),
            .in2(N__24197),
            .in3(N__23588),
            .lcout(\QuadInstance1.Quad_RNIPI0OZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNIQJ0O_3_LC_14_6_7 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_RNIQJ0O_3_LC_14_6_7 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNIQJ0O_3_LC_14_6_7 .LUT_INIT=16'b1010111100000000;
    LogicCell40 \QuadInstance1.Quad_RNIQJ0O_3_LC_14_6_7  (
            .in0(N__24006),
            .in1(N__27878),
            .in2(N__23611),
            .in3(N__24173),
            .lcout(\QuadInstance1.Quad_RNIQJ0OZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNIAR5D_12_LC_14_7_0 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_RNIAR5D_12_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNIAR5D_12_LC_14_7_0 .LUT_INIT=16'b1010101000100010;
    LogicCell40 \QuadInstance1.Quad_RNIAR5D_12_LC_14_7_0  (
            .in0(N__24200),
            .in1(N__23618),
            .in2(N__24128),
            .in3(N__24022),
            .lcout(\QuadInstance1.Quad_RNIAR5DZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNIBS5D_13_LC_14_7_1 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_RNIBS5D_13_LC_14_7_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNIBS5D_13_LC_14_7_1 .LUT_INIT=16'b1000110010001100;
    LogicCell40 \QuadInstance1.Quad_RNIBS5D_13_LC_14_7_1  (
            .in0(N__24023),
            .in1(N__24201),
            .in2(N__23625),
            .in3(N__23918),
            .lcout(\QuadInstance1.Quad_RNIBS5DZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNICT5D_14_LC_14_7_2 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_RNICT5D_14_LC_14_7_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNICT5D_14_LC_14_7_2 .LUT_INIT=16'b1111000000110000;
    LogicCell40 \QuadInstance1.Quad_RNICT5D_14_LC_14_7_2  (
            .in0(N__28190),
            .in1(N__23622),
            .in2(N__24209),
            .in3(N__24024),
            .lcout(\QuadInstance1.Quad_RNICT5DZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNIVO0O_8_LC_14_7_3 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_RNIVO0O_8_LC_14_7_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNIVO0O_8_LC_14_7_3 .LUT_INIT=16'b1010111100000000;
    LogicCell40 \QuadInstance1.Quad_RNIVO0O_8_LC_14_7_3  (
            .in0(N__24021),
            .in1(N__37013),
            .in2(N__23624),
            .in3(N__24199),
            .lcout(\QuadInstance1.Quad_RNIVO0OZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_RNO_0_15_LC_14_7_4 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_RNO_0_15_LC_14_7_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance1.Quad_RNO_0_15_LC_14_7_4 .LUT_INIT=16'b0101101010011010;
    LogicCell40 \QuadInstance1.Quad_RNO_0_15_LC_14_7_4  (
            .in0(N__24227),
            .in1(N__23623),
            .in2(N__24210),
            .in3(N__24025),
            .lcout(\QuadInstance1.un1_Quad_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.Quad_0_LC_14_7_5 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_0_LC_14_7_5 .SEQ_MODE=4'b1000;
    defparam \QuadInstance1.Quad_0_LC_14_7_5 .LUT_INIT=16'b1000110111011000;
    LogicCell40 \QuadInstance1.Quad_0_LC_14_7_5  (
            .in0(N__24027),
            .in1(N__31411),
            .in2(N__30947),
            .in3(N__24208),
            .lcout(dataRead1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38674),
            .ce(),
            .sr(N__35734));
    defparam \QuadInstance1.Quad_12_LC_14_7_6 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_12_LC_14_7_6 .SEQ_MODE=4'b1000;
    defparam \QuadInstance1.Quad_12_LC_14_7_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance1.Quad_12_LC_14_7_6  (
            .in0(N__28833),
            .in1(N__24028),
            .in2(_gnd_net_),
            .in3(N__24135),
            .lcout(dataRead1_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38674),
            .ce(),
            .sr(N__35734));
    defparam \QuadInstance1.Quad_13_LC_14_7_7 .C_ON=1'b0;
    defparam \QuadInstance1.Quad_13_LC_14_7_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance1.Quad_13_LC_14_7_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance1.Quad_13_LC_14_7_7  (
            .in0(N__24026),
            .in1(N__28715),
            .in2(_gnd_net_),
            .in3(N__23928),
            .lcout(dataRead1_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38674),
            .ce(),
            .sr(N__35734));
    defparam OutReg_ess_RNO_2_1_LC_14_8_0.C_ON=1'b0;
    defparam OutReg_ess_RNO_2_1_LC_14_8_0.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_2_1_LC_14_8_0.LUT_INIT=16'b1011100000110011;
    LogicCell40 OutReg_ess_RNO_2_1_LC_14_8_0 (
            .in0(N__23897),
            .in1(N__23751),
            .in2(N__23868),
            .in3(N__32926),
            .lcout(),
            .ltout(OutReg_ess_RNO_2Z0Z_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_0_1_LC_14_8_1.C_ON=1'b0;
    defparam OutReg_ess_RNO_0_1_LC_14_8_1.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_0_1_LC_14_8_1.LUT_INIT=16'b1111110000110000;
    LogicCell40 OutReg_ess_RNO_0_1_LC_14_8_1 (
            .in0(_gnd_net_),
            .in1(N__37502),
            .in2(N__23838),
            .in3(N__23757),
            .lcout(OutReg_ess_RNO_0Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_3_1_LC_14_8_2.C_ON=1'b0;
    defparam OutReg_ess_RNO_3_1_LC_14_8_2.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_3_1_LC_14_8_2.LUT_INIT=16'b0011000100111101;
    LogicCell40 OutReg_ess_RNO_3_1_LC_14_8_2 (
            .in0(N__23827),
            .in1(N__34732),
            .in2(N__34884),
            .in3(N__23800),
            .lcout(),
            .ltout(OutReg_0_4_i_m3_ns_1_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_1_1_LC_14_8_3.C_ON=1'b0;
    defparam OutReg_ess_RNO_1_1_LC_14_8_3.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_1_1_LC_14_8_3.LUT_INIT=16'b1100101000001111;
    LogicCell40 OutReg_ess_RNO_1_1_LC_14_8_3 (
            .in0(N__25834),
            .in1(N__23787),
            .in2(N__23760),
            .in3(N__32811),
            .lcout(OutReg_ess_RNO_1Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_4_1_LC_14_8_4.C_ON=1'b0;
    defparam OutReg_ess_RNO_4_1_LC_14_8_4.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_4_1_LC_14_8_4.LUT_INIT=16'b0011000100111101;
    LogicCell40 OutReg_ess_RNO_4_1_LC_14_8_4 (
            .in0(N__32716),
            .in1(N__28102),
            .in2(N__27996),
            .in3(N__27220),
            .lcout(OutReg_0_5_i_m3_ns_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_received_fast_esr_2_LC_14_8_5.C_ON=1'b0;
    defparam data_received_fast_esr_2_LC_14_8_5.SEQ_MODE=4'b1000;
    defparam data_received_fast_esr_2_LC_14_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 data_received_fast_esr_2_LC_14_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37504),
            .lcout(data_received_fastZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38665),
            .ce(N__26178),
            .sr(N__26156));
    defparam data_received_2_rep1_esr_LC_14_8_6.C_ON=1'b0;
    defparam data_received_2_rep1_esr_LC_14_8_6.SEQ_MODE=4'b1000;
    defparam data_received_2_rep1_esr_LC_14_8_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 data_received_2_rep1_esr_LC_14_8_6 (
            .in0(N__37503),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(data_received_2_repZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38665),
            .ce(N__26178),
            .sr(N__26156));
    defparam OutReg_ess_RNO_3_3_LC_14_8_7.C_ON=1'b0;
    defparam OutReg_ess_RNO_3_3_LC_14_8_7.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_3_3_LC_14_8_7.LUT_INIT=16'b0101010100011011;
    LogicCell40 OutReg_ess_RNO_3_3_LC_14_8_7 (
            .in0(N__34733),
            .in1(N__24410),
            .in2(N__24374),
            .in3(N__34862),
            .lcout(OutReg_0_4_i_m3_ns_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_15_LC_14_9_0.C_ON=1'b0;
    defparam OutReg_ess_15_LC_14_9_0.SEQ_MODE=4'b1001;
    defparam OutReg_ess_15_LC_14_9_0.LUT_INIT=16'b1111000111100000;
    LogicCell40 OutReg_ess_15_LC_14_9_0 (
            .in0(N__38946),
            .in1(N__37374),
            .in2(N__26205),
            .in3(N__37821),
            .lcout(OutRegZ0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38653),
            .ce(N__37245),
            .sr(N__37135));
    defparam OutReg_ess_RNO_3_15_LC_14_9_1.C_ON=1'b0;
    defparam OutReg_ess_RNO_3_15_LC_14_9_1.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_3_15_LC_14_9_1.LUT_INIT=16'b0000111101010011;
    LogicCell40 OutReg_ess_RNO_3_15_LC_14_9_1 (
            .in0(N__24336),
            .in1(N__24315),
            .in2(N__28016),
            .in3(N__28101),
            .lcout(),
            .ltout(OutReg_0_4_i_m3_ns_1_15_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_1_15_LC_14_9_2.C_ON=1'b0;
    defparam OutReg_ess_RNO_1_15_LC_14_9_2.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_1_15_LC_14_9_2.LUT_INIT=16'b1100101000001111;
    LogicCell40 OutReg_ess_RNO_1_15_LC_14_9_2 (
            .in0(N__24291),
            .in1(N__24269),
            .in2(N__24249),
            .in3(N__37708),
            .lcout(OutReg_ess_RNO_1Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_2_15_LC_14_9_4.C_ON=1'b0;
    defparam OutReg_ess_RNO_2_15_LC_14_9_4.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_2_15_LC_14_9_4.LUT_INIT=16'b1110010001010101;
    LogicCell40 OutReg_ess_RNO_2_15_LC_14_9_4 (
            .in0(N__25197),
            .in1(N__24246),
            .in2(N__24228),
            .in3(N__38114),
            .lcout(OutReg_ess_RNO_2Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_received_esr_5_LC_14_10_1.C_ON=1'b0;
    defparam data_received_esr_5_LC_14_10_1.SEQ_MODE=4'b1000;
    defparam data_received_esr_5_LC_14_10_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 data_received_esr_5_LC_14_10_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34979),
            .lcout(data_receivedZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38643),
            .ce(N__26183),
            .sr(N__26153));
    defparam data_received_esr_7_LC_14_10_2.C_ON=1'b0;
    defparam data_received_esr_7_LC_14_10_2.SEQ_MODE=4'b1000;
    defparam data_received_esr_7_LC_14_10_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 data_received_esr_7_LC_14_10_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24437),
            .lcout(data_receivedZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38643),
            .ce(N__26183),
            .sr(N__26153));
    defparam data_received_esr_9_LC_14_10_4.C_ON=1'b0;
    defparam data_received_esr_9_LC_14_10_4.SEQ_MODE=4'b1000;
    defparam data_received_esr_9_LC_14_10_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 data_received_esr_9_LC_14_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24485),
            .lcout(data_receivedZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38643),
            .ce(N__26183),
            .sr(N__26153));
    defparam data_received_esr_22_LC_14_10_5.C_ON=1'b0;
    defparam data_received_esr_22_LC_14_10_5.SEQ_MODE=4'b1000;
    defparam data_received_esr_22_LC_14_10_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 data_received_esr_22_LC_14_10_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33842),
            .lcout(data_receivedZ0Z_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38643),
            .ce(N__26183),
            .sr(N__26153));
    defparam data_received_esr_6_LC_14_10_6.C_ON=1'b0;
    defparam data_received_esr_6_LC_14_10_6.SEQ_MODE=4'b1000;
    defparam data_received_esr_6_LC_14_10_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 data_received_esr_6_LC_14_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24449),
            .lcout(data_receivedZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38643),
            .ce(N__26183),
            .sr(N__26153));
    defparam data_received_esr_8_LC_14_10_7.C_ON=1'b0;
    defparam data_received_esr_8_LC_14_10_7.SEQ_MODE=4'b1000;
    defparam data_received_esr_8_LC_14_10_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 data_received_esr_8_LC_14_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24425),
            .lcout(data_receivedZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38643),
            .ce(N__26183),
            .sr(N__26153));
    defparam dataWrite_2_LC_14_11_0.C_ON=1'b0;
    defparam dataWrite_2_LC_14_11_0.SEQ_MODE=4'b1000;
    defparam dataWrite_2_LC_14_11_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 dataWrite_2_LC_14_11_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37712),
            .lcout(dataWriteZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38634),
            .ce(N__24462),
            .sr(_gnd_net_));
    defparam dataWrite_3_LC_14_11_1.C_ON=1'b0;
    defparam dataWrite_3_LC_14_11_1.SEQ_MODE=4'b1000;
    defparam dataWrite_3_LC_14_11_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 dataWrite_3_LC_14_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30638),
            .lcout(dataWriteZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38634),
            .ce(N__24462),
            .sr(_gnd_net_));
    defparam dataWrite_4_LC_14_11_2.C_ON=1'b0;
    defparam dataWrite_4_LC_14_11_2.SEQ_MODE=4'b1000;
    defparam dataWrite_4_LC_14_11_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 dataWrite_4_LC_14_11_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34978),
            .lcout(dataWriteZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38634),
            .ce(N__24462),
            .sr(_gnd_net_));
    defparam dataWrite_5_LC_14_11_3.C_ON=1'b0;
    defparam dataWrite_5_LC_14_11_3.SEQ_MODE=4'b1000;
    defparam dataWrite_5_LC_14_11_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 dataWrite_5_LC_14_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24450),
            .lcout(dataWriteZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38634),
            .ce(N__24462),
            .sr(_gnd_net_));
    defparam dataWrite_6_LC_14_11_4.C_ON=1'b0;
    defparam dataWrite_6_LC_14_11_4.SEQ_MODE=4'b1000;
    defparam dataWrite_6_LC_14_11_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 dataWrite_6_LC_14_11_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24438),
            .lcout(dataWriteZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38634),
            .ce(N__24462),
            .sr(_gnd_net_));
    defparam dataWrite_7_LC_14_11_5.C_ON=1'b0;
    defparam dataWrite_7_LC_14_11_5.SEQ_MODE=4'b1000;
    defparam dataWrite_7_LC_14_11_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 dataWrite_7_LC_14_11_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24426),
            .lcout(dataWriteZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38634),
            .ce(N__24462),
            .sr(_gnd_net_));
    defparam dataWrite_8_LC_14_11_6.C_ON=1'b0;
    defparam dataWrite_8_LC_14_11_6.SEQ_MODE=4'b1000;
    defparam dataWrite_8_LC_14_11_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 dataWrite_8_LC_14_11_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24486),
            .lcout(dataWriteZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38634),
            .ce(N__24462),
            .sr(_gnd_net_));
    defparam dataWrite_9_LC_14_11_7.C_ON=1'b0;
    defparam dataWrite_9_LC_14_11_7.SEQ_MODE=4'b1000;
    defparam dataWrite_9_LC_14_11_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 dataWrite_9_LC_14_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24473),
            .lcout(dataWriteZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38634),
            .ce(N__24462),
            .sr(_gnd_net_));
    defparam \PWMInstance3.PWMPulseWidthCount_esr_11_LC_14_12_0 .C_ON=1'b0;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_11_LC_14_12_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_11_LC_14_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance3.PWMPulseWidthCount_esr_11_LC_14_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35974),
            .lcout(\PWMInstance3.PWMPulseWidthCountZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38621),
            .ce(N__29290),
            .sr(N__35765));
    defparam \PWMInstance3.PWMPulseWidthCount_esr_8_LC_14_12_2 .C_ON=1'b0;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_8_LC_14_12_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_8_LC_14_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance3.PWMPulseWidthCount_esr_8_LC_14_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28912),
            .lcout(\PWMInstance3.PWMPulseWidthCountZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38621),
            .ce(N__29290),
            .sr(N__35765));
    defparam \PWMInstance3.PWMPulseWidthCount_esr_5_LC_14_12_3 .C_ON=1'b0;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_5_LC_14_12_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_5_LC_14_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance3.PWMPulseWidthCount_esr_5_LC_14_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36284),
            .lcout(\PWMInstance3.PWMPulseWidthCountZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38621),
            .ce(N__29290),
            .sr(N__35765));
    defparam \PWMInstance3.PWMPulseWidthCount_esr_10_LC_14_12_4 .C_ON=1'b0;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_10_LC_14_12_4 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_10_LC_14_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance3.PWMPulseWidthCount_esr_10_LC_14_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36157),
            .lcout(\PWMInstance3.PWMPulseWidthCountZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38621),
            .ce(N__29290),
            .sr(N__35765));
    defparam \PWMInstance3.PWMPulseWidthCount_esr_3_LC_14_12_6 .C_ON=1'b0;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_3_LC_14_12_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_3_LC_14_12_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \PWMInstance3.PWMPulseWidthCount_esr_3_LC_14_12_6  (
            .in0(_gnd_net_),
            .in1(N__31985),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PWMInstance3.PWMPulseWidthCountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38621),
            .ce(N__29290),
            .sr(N__35765));
    defparam \PWMInstance3.out_RNO_0_LC_14_13_0 .C_ON=1'b0;
    defparam \PWMInstance3.out_RNO_0_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance3.out_RNO_0_LC_14_13_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \PWMInstance3.out_RNO_0_LC_14_13_0  (
            .in0(N__24621),
            .in1(N__24604),
            .in2(N__26709),
            .in3(N__24589),
            .lcout(\PWMInstance3.un1_periodCounter12_1_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance3.clkCount_0_LC_14_13_1 .C_ON=1'b0;
    defparam \PWMInstance3.clkCount_0_LC_14_13_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.clkCount_0_LC_14_13_1 .LUT_INIT=16'b1010101000000101;
    LogicCell40 \PWMInstance3.clkCount_0_LC_14_13_1  (
            .in0(N__24590),
            .in1(_gnd_net_),
            .in2(N__24611),
            .in3(N__24635),
            .lcout(\PWMInstance3.clkCountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38612),
            .ce(),
            .sr(N__35771));
    defparam \PWMInstance3.PWMPulseWidthCount_esr_ctle_15_LC_14_13_2 .C_ON=1'b0;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_ctle_15_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_ctle_15_LC_14_13_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \PWMInstance3.PWMPulseWidthCount_esr_ctle_15_LC_14_13_2  (
            .in0(N__35830),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24634),
            .lcout(\PWMInstance3.pwmWrite_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance3.clkCount_1_LC_14_13_3 .C_ON=1'b0;
    defparam \PWMInstance3.clkCount_1_LC_14_13_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.clkCount_1_LC_14_13_3 .LUT_INIT=16'b1111000000001010;
    LogicCell40 \PWMInstance3.clkCount_1_LC_14_13_3  (
            .in0(N__24591),
            .in1(_gnd_net_),
            .in2(N__24612),
            .in3(N__24636),
            .lcout(\PWMInstance3.clkCountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38612),
            .ce(),
            .sr(N__35771));
    defparam \PWMInstance3.clkCount_RNI21FG_0_LC_14_13_4 .C_ON=1'b0;
    defparam \PWMInstance3.clkCount_RNI21FG_0_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance3.clkCount_RNI21FG_0_LC_14_13_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \PWMInstance3.clkCount_RNI21FG_0_LC_14_13_4  (
            .in0(N__24620),
            .in1(N__24603),
            .in2(_gnd_net_),
            .in3(N__24588),
            .lcout(\PWMInstance3.periodCounter12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance3.periodCounter_RNI8K3C_16_LC_14_13_5 .C_ON=1'b0;
    defparam \PWMInstance3.periodCounter_RNI8K3C_16_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \PWMInstance3.periodCounter_RNI8K3C_16_LC_14_13_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \PWMInstance3.periodCounter_RNI8K3C_16_LC_14_13_5  (
            .in0(_gnd_net_),
            .in1(N__26705),
            .in2(_gnd_net_),
            .in3(N__29497),
            .lcout(),
            .ltout(\PWMInstance3.un1_periodCounter12_1_0_a2_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance3.periodCounter_RNIB2M81_1_LC_14_13_6 .C_ON=1'b0;
    defparam \PWMInstance3.periodCounter_RNIB2M81_1_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \PWMInstance3.periodCounter_RNIB2M81_1_LC_14_13_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \PWMInstance3.periodCounter_RNIB2M81_1_LC_14_13_6  (
            .in0(N__29038),
            .in1(N__29170),
            .in2(N__24576),
            .in3(N__26428),
            .lcout(),
            .ltout(\PWMInstance3.un1_periodCounter12_1_0_a2_0_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance3.periodCounter_RNI0E0J3_0_LC_14_13_7 .C_ON=1'b0;
    defparam \PWMInstance3.periodCounter_RNI0E0J3_0_LC_14_13_7 .SEQ_MODE=4'b0000;
    defparam \PWMInstance3.periodCounter_RNI0E0J3_0_LC_14_13_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \PWMInstance3.periodCounter_RNI0E0J3_0_LC_14_13_7  (
            .in0(N__28389),
            .in1(N__29067),
            .in2(N__24573),
            .in3(N__26457),
            .lcout(\PWMInstance3.out_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance6.PWMPulseWidthCount_esr_9_LC_14_14_4 .C_ON=1'b0;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_9_LC_14_14_4 .SEQ_MODE=4'b1000;
    defparam \PWMInstance6.PWMPulseWidthCount_esr_9_LC_14_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance6.PWMPulseWidthCount_esr_9_LC_14_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28523),
            .lcout(\PWMInstance6.PWMPulseWidthCountZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38600),
            .ce(N__24552),
            .sr(N__35775));
    defparam \PWMInstance4.periodCounter_RNIRPSE_3_LC_14_15_0 .C_ON=1'b0;
    defparam \PWMInstance4.periodCounter_RNIRPSE_3_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance4.periodCounter_RNIRPSE_3_LC_14_15_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \PWMInstance4.periodCounter_RNIRPSE_3_LC_14_15_0  (
            .in0(N__26550),
            .in1(N__24832),
            .in2(N__24780),
            .in3(N__24673),
            .lcout(\PWMInstance4.un1_periodCounter12_1_0_a2_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_14_15_1 .C_ON=1'b0;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_14_15_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_14_15_1 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance4.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_14_15_1  (
            .in0(N__24498),
            .in1(N__24492),
            .in2(N__24675),
            .in3(N__24695),
            .lcout(\PWMInstance4.un1_PWMPulseWidthCount_0_I_9_c_RNO_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance4.PWMPulseWidthCount_esr_2_LC_14_15_2 .C_ON=1'b0;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_2_LC_14_15_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_2_LC_14_15_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \PWMInstance4.PWMPulseWidthCount_esr_2_LC_14_15_2  (
            .in0(N__31543),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PWMInstance4.PWMPulseWidthCountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38593),
            .ce(N__26954),
            .sr(N__35783));
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_14_15_4 .C_ON=1'b0;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_14_15_4 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance4.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_14_15_4  (
            .in0(N__24717),
            .in1(N__24723),
            .in2(N__26841),
            .in3(N__24915),
            .lcout(\PWMInstance4.un1_PWMPulseWidthCount_0_I_21_c_RNO_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance4.PWMPulseWidthCount_esr_14_LC_14_15_5 .C_ON=1'b0;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_14_LC_14_15_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_14_LC_14_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance4.PWMPulseWidthCount_esr_14_LC_14_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34395),
            .lcout(\PWMInstance4.PWMPulseWidthCountZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38593),
            .ce(N__26954),
            .sr(N__35783));
    defparam \PWMInstance4.PWMPulseWidthCount_esr_15_LC_14_15_6 .C_ON=1'b0;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_15_LC_14_15_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_15_LC_14_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance4.PWMPulseWidthCount_esr_15_LC_14_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31858),
            .lcout(\PWMInstance4.PWMPulseWidthCountZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38593),
            .ce(N__26954),
            .sr(N__35783));
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_14_15_7 .C_ON=1'b0;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_14_15_7 .SEQ_MODE=4'b0000;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_14_15_7 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \PWMInstance4.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_14_15_7  (
            .in0(N__24711),
            .in1(N__24705),
            .in2(N__26688),
            .in3(N__24750),
            .lcout(\PWMInstance4.un1_PWMPulseWidthCount_0_I_39_c_RNO_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance4.periodCounter_0_LC_14_16_0 .C_ON=1'b1;
    defparam \PWMInstance4.periodCounter_0_LC_14_16_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.periodCounter_0_LC_14_16_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance4.periodCounter_0_LC_14_16_0  (
            .in0(_gnd_net_),
            .in1(N__26664),
            .in2(N__26856),
            .in3(N__26855),
            .lcout(\PWMInstance4.periodCounterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_14_16_0_),
            .carryout(\PWMInstance4.un1_periodCounter_2_cry_0 ),
            .clk(N__38582),
            .ce(),
            .sr(N__35297));
    defparam \PWMInstance4.periodCounter_1_LC_14_16_1 .C_ON=1'b1;
    defparam \PWMInstance4.periodCounter_1_LC_14_16_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.periodCounter_1_LC_14_16_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance4.periodCounter_1_LC_14_16_1  (
            .in0(_gnd_net_),
            .in1(N__26813),
            .in2(_gnd_net_),
            .in3(N__24699),
            .lcout(\PWMInstance4.periodCounterZ0Z_1 ),
            .ltout(),
            .carryin(\PWMInstance4.un1_periodCounter_2_cry_0 ),
            .carryout(\PWMInstance4.un1_periodCounter_2_cry_1 ),
            .clk(N__38582),
            .ce(),
            .sr(N__35297));
    defparam \PWMInstance4.periodCounter_2_LC_14_16_2 .C_ON=1'b1;
    defparam \PWMInstance4.periodCounter_2_LC_14_16_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.periodCounter_2_LC_14_16_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance4.periodCounter_2_LC_14_16_2  (
            .in0(_gnd_net_),
            .in1(N__24696),
            .in2(_gnd_net_),
            .in3(N__24678),
            .lcout(\PWMInstance4.periodCounterZ0Z_2 ),
            .ltout(),
            .carryin(\PWMInstance4.un1_periodCounter_2_cry_1 ),
            .carryout(\PWMInstance4.un1_periodCounter_2_cry_2 ),
            .clk(N__38582),
            .ce(),
            .sr(N__35297));
    defparam \PWMInstance4.periodCounter_3_LC_14_16_3 .C_ON=1'b1;
    defparam \PWMInstance4.periodCounter_3_LC_14_16_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.periodCounter_3_LC_14_16_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance4.periodCounter_3_LC_14_16_3  (
            .in0(_gnd_net_),
            .in1(N__24674),
            .in2(_gnd_net_),
            .in3(N__24657),
            .lcout(\PWMInstance4.periodCounterZ0Z_3 ),
            .ltout(),
            .carryin(\PWMInstance4.un1_periodCounter_2_cry_2 ),
            .carryout(\PWMInstance4.un1_periodCounter_2_cry_3 ),
            .clk(N__38582),
            .ce(),
            .sr(N__35297));
    defparam \PWMInstance4.periodCounter_4_LC_14_16_4 .C_ON=1'b1;
    defparam \PWMInstance4.periodCounter_4_LC_14_16_4 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.periodCounter_4_LC_14_16_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance4.periodCounter_4_LC_14_16_4  (
            .in0(_gnd_net_),
            .in1(N__24654),
            .in2(_gnd_net_),
            .in3(N__24639),
            .lcout(\PWMInstance4.periodCounterZ0Z_4 ),
            .ltout(),
            .carryin(\PWMInstance4.un1_periodCounter_2_cry_3 ),
            .carryout(\PWMInstance4.un1_periodCounter_2_cry_4 ),
            .clk(N__38582),
            .ce(),
            .sr(N__35297));
    defparam \PWMInstance4.periodCounter_5_LC_14_16_5 .C_ON=1'b1;
    defparam \PWMInstance4.periodCounter_5_LC_14_16_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.periodCounter_5_LC_14_16_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance4.periodCounter_5_LC_14_16_5  (
            .in0(_gnd_net_),
            .in1(N__24833),
            .in2(_gnd_net_),
            .in3(N__24813),
            .lcout(\PWMInstance4.periodCounterZ0Z_5 ),
            .ltout(),
            .carryin(\PWMInstance4.un1_periodCounter_2_cry_4 ),
            .carryout(\PWMInstance4.un1_periodCounter_2_cry_5 ),
            .clk(N__38582),
            .ce(),
            .sr(N__35297));
    defparam \PWMInstance4.periodCounter_6_LC_14_16_6 .C_ON=1'b1;
    defparam \PWMInstance4.periodCounter_6_LC_14_16_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.periodCounter_6_LC_14_16_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance4.periodCounter_6_LC_14_16_6  (
            .in0(_gnd_net_),
            .in1(N__26619),
            .in2(_gnd_net_),
            .in3(N__24810),
            .lcout(\PWMInstance4.periodCounterZ0Z_6 ),
            .ltout(),
            .carryin(\PWMInstance4.un1_periodCounter_2_cry_5 ),
            .carryout(\PWMInstance4.un1_periodCounter_2_cry_6 ),
            .clk(N__38582),
            .ce(),
            .sr(N__35297));
    defparam \PWMInstance4.periodCounter_7_LC_14_16_7 .C_ON=1'b1;
    defparam \PWMInstance4.periodCounter_7_LC_14_16_7 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.periodCounter_7_LC_14_16_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance4.periodCounter_7_LC_14_16_7  (
            .in0(N__26749),
            .in1(N__26994),
            .in2(_gnd_net_),
            .in3(N__24807),
            .lcout(\PWMInstance4.periodCounterZ0Z_7 ),
            .ltout(),
            .carryin(\PWMInstance4.un1_periodCounter_2_cry_6 ),
            .carryout(\PWMInstance4.un1_periodCounter_2_cry_7 ),
            .clk(N__38582),
            .ce(),
            .sr(N__35297));
    defparam \PWMInstance4.periodCounter_8_LC_14_17_0 .C_ON=1'b1;
    defparam \PWMInstance4.periodCounter_8_LC_14_17_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.periodCounter_8_LC_14_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance4.periodCounter_8_LC_14_17_0  (
            .in0(_gnd_net_),
            .in1(N__26567),
            .in2(_gnd_net_),
            .in3(N__24804),
            .lcout(\PWMInstance4.periodCounterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_14_17_0_),
            .carryout(\PWMInstance4.un1_periodCounter_2_cry_8 ),
            .clk(N__38572),
            .ce(),
            .sr(N__35295));
    defparam \PWMInstance4.periodCounter_9_LC_14_17_1 .C_ON=1'b1;
    defparam \PWMInstance4.periodCounter_9_LC_14_17_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.periodCounter_9_LC_14_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance4.periodCounter_9_LC_14_17_1  (
            .in0(_gnd_net_),
            .in1(N__26548),
            .in2(_gnd_net_),
            .in3(N__24801),
            .lcout(\PWMInstance4.periodCounterZ0Z_9 ),
            .ltout(),
            .carryin(\PWMInstance4.un1_periodCounter_2_cry_8 ),
            .carryout(\PWMInstance4.un1_periodCounter_2_cry_9 ),
            .clk(N__38572),
            .ce(),
            .sr(N__35295));
    defparam \PWMInstance4.periodCounter_10_LC_14_17_2 .C_ON=1'b1;
    defparam \PWMInstance4.periodCounter_10_LC_14_17_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.periodCounter_10_LC_14_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance4.periodCounter_10_LC_14_17_2  (
            .in0(_gnd_net_),
            .in1(N__24798),
            .in2(_gnd_net_),
            .in3(N__24783),
            .lcout(\PWMInstance4.periodCounterZ0Z_10 ),
            .ltout(),
            .carryin(\PWMInstance4.un1_periodCounter_2_cry_9 ),
            .carryout(\PWMInstance4.un1_periodCounter_2_cry_10 ),
            .clk(N__38572),
            .ce(),
            .sr(N__35295));
    defparam \PWMInstance4.periodCounter_11_LC_14_17_3 .C_ON=1'b1;
    defparam \PWMInstance4.periodCounter_11_LC_14_17_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.periodCounter_11_LC_14_17_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance4.periodCounter_11_LC_14_17_3  (
            .in0(N__26747),
            .in1(N__24775),
            .in2(_gnd_net_),
            .in3(N__24753),
            .lcout(\PWMInstance4.periodCounterZ0Z_11 ),
            .ltout(),
            .carryin(\PWMInstance4.un1_periodCounter_2_cry_10 ),
            .carryout(\PWMInstance4.un1_periodCounter_2_cry_11 ),
            .clk(N__38572),
            .ce(),
            .sr(N__35295));
    defparam \PWMInstance4.periodCounter_12_LC_14_17_4 .C_ON=1'b1;
    defparam \PWMInstance4.periodCounter_12_LC_14_17_4 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.periodCounter_12_LC_14_17_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance4.periodCounter_12_LC_14_17_4  (
            .in0(N__26746),
            .in1(N__24749),
            .in2(_gnd_net_),
            .in3(N__24729),
            .lcout(\PWMInstance4.periodCounterZ0Z_12 ),
            .ltout(),
            .carryin(\PWMInstance4.un1_periodCounter_2_cry_11 ),
            .carryout(\PWMInstance4.un1_periodCounter_2_cry_12 ),
            .clk(N__38572),
            .ce(),
            .sr(N__35295));
    defparam \PWMInstance4.periodCounter_13_LC_14_17_5 .C_ON=1'b1;
    defparam \PWMInstance4.periodCounter_13_LC_14_17_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.periodCounter_13_LC_14_17_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance4.periodCounter_13_LC_14_17_5  (
            .in0(N__26748),
            .in1(N__26683),
            .in2(_gnd_net_),
            .in3(N__24726),
            .lcout(\PWMInstance4.periodCounterZ0Z_13 ),
            .ltout(),
            .carryin(\PWMInstance4.un1_periodCounter_2_cry_12 ),
            .carryout(\PWMInstance4.un1_periodCounter_2_cry_13 ),
            .clk(N__38572),
            .ce(),
            .sr(N__35295));
    defparam \PWMInstance4.periodCounter_14_LC_14_17_6 .C_ON=1'b1;
    defparam \PWMInstance4.periodCounter_14_LC_14_17_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.periodCounter_14_LC_14_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance4.periodCounter_14_LC_14_17_6  (
            .in0(_gnd_net_),
            .in1(N__24914),
            .in2(_gnd_net_),
            .in3(N__24894),
            .lcout(\PWMInstance4.periodCounterZ0Z_14 ),
            .ltout(),
            .carryin(\PWMInstance4.un1_periodCounter_2_cry_13 ),
            .carryout(\PWMInstance4.un1_periodCounter_2_cry_14 ),
            .clk(N__38572),
            .ce(),
            .sr(N__35295));
    defparam \PWMInstance4.periodCounter_15_LC_14_17_7 .C_ON=1'b1;
    defparam \PWMInstance4.periodCounter_15_LC_14_17_7 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.periodCounter_15_LC_14_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance4.periodCounter_15_LC_14_17_7  (
            .in0(_gnd_net_),
            .in1(N__26834),
            .in2(_gnd_net_),
            .in3(N__24891),
            .lcout(\PWMInstance4.periodCounterZ0Z_15 ),
            .ltout(),
            .carryin(\PWMInstance4.un1_periodCounter_2_cry_14 ),
            .carryout(\PWMInstance4.un1_periodCounter_2_cry_15 ),
            .clk(N__38572),
            .ce(),
            .sr(N__35295));
    defparam \PWMInstance4.periodCounter_16_LC_14_18_0 .C_ON=1'b0;
    defparam \PWMInstance4.periodCounter_16_LC_14_18_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.periodCounter_16_LC_14_18_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance4.periodCounter_16_LC_14_18_0  (
            .in0(N__26750),
            .in1(N__27009),
            .in2(_gnd_net_),
            .in3(N__24888),
            .lcout(\PWMInstance4.periodCounterZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38564),
            .ce(),
            .sr(N__35293));
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_1_c_LC_15_1_0 .C_ON=1'b1;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_1_c_LC_15_1_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_1_c_LC_15_1_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance4.un1_PWMPulseWidthCount_0_I_1_c_LC_15_1_0  (
            .in0(_gnd_net_),
            .in1(N__26637),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_1_0_),
            .carryout(\PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_9_c_LC_15_1_1 .C_ON=1'b1;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_9_c_LC_15_1_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_9_c_LC_15_1_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance4.un1_PWMPulseWidthCount_0_I_9_c_LC_15_1_1  (
            .in0(_gnd_net_),
            .in1(N__24885),
            .in2(N__32544),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_0 ),
            .carryout(\PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_15_c_LC_15_1_2 .C_ON=1'b1;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_15_c_LC_15_1_2 .SEQ_MODE=4'b0000;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_15_c_LC_15_1_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance4.un1_PWMPulseWidthCount_0_I_15_c_LC_15_1_2  (
            .in0(_gnd_net_),
            .in1(N__24867),
            .in2(N__32538),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_1 ),
            .carryout(\PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_27_c_LC_15_1_3 .C_ON=1'b1;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_27_c_LC_15_1_3 .SEQ_MODE=4'b0000;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_27_c_LC_15_1_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance4.un1_PWMPulseWidthCount_0_I_27_c_LC_15_1_3  (
            .in0(_gnd_net_),
            .in1(N__26604),
            .in2(N__32542),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_2 ),
            .carryout(\PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_45_c_LC_15_1_4 .C_ON=1'b1;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_45_c_LC_15_1_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_45_c_LC_15_1_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance4.un1_PWMPulseWidthCount_0_I_45_c_LC_15_1_4  (
            .in0(_gnd_net_),
            .in1(N__26517),
            .in2(N__32540),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_3 ),
            .carryout(\PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_33_c_LC_15_1_5 .C_ON=1'b1;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_33_c_LC_15_1_5 .SEQ_MODE=4'b0000;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_33_c_LC_15_1_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance4.un1_PWMPulseWidthCount_0_I_33_c_LC_15_1_5  (
            .in0(_gnd_net_),
            .in1(N__24852),
            .in2(N__32543),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_4 ),
            .carryout(\PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_39_c_LC_15_1_6 .C_ON=1'b1;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_39_c_LC_15_1_6 .SEQ_MODE=4'b0000;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_39_c_LC_15_1_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance4.un1_PWMPulseWidthCount_0_I_39_c_LC_15_1_6  (
            .in0(_gnd_net_),
            .in1(N__25020),
            .in2(N__32539),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_5 ),
            .carryout(\PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_21_c_LC_15_1_7 .C_ON=1'b1;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_21_c_LC_15_1_7 .SEQ_MODE=4'b0000;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_21_c_LC_15_1_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance4.un1_PWMPulseWidthCount_0_I_21_c_LC_15_1_7  (
            .in0(_gnd_net_),
            .in1(N__25002),
            .in2(N__32541),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_6 ),
            .carryout(\PWMInstance4.un1_PWMPulseWidthCount_0_data_tmp_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance4.out_LC_15_2_0 .C_ON=1'b0;
    defparam \PWMInstance4.out_LC_15_2_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.out_LC_15_2_0 .LUT_INIT=16'b1111101011110010;
    LogicCell40 \PWMInstance4.out_LC_15_2_0  (
            .in0(N__24962),
            .in1(N__27021),
            .in2(N__26757),
            .in3(N__24984),
            .lcout(PWM4_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38717),
            .ce(),
            .sr(N__35701));
    defparam \QuadInstance4.un1_Quad_cry_0_c_LC_15_3_0 .C_ON=1'b1;
    defparam \QuadInstance4.un1_Quad_cry_0_c_LC_15_3_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.un1_Quad_cry_0_c_LC_15_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \QuadInstance4.un1_Quad_cry_0_c_LC_15_3_0  (
            .in0(_gnd_net_),
            .in1(N__27432),
            .in2(N__30284),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_3_0_),
            .carryout(\QuadInstance4.un1_Quad_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_RNO_0_1_LC_15_3_1 .C_ON=1'b1;
    defparam \QuadInstance4.Quad_RNO_0_1_LC_15_3_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNO_0_1_LC_15_3_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance4.Quad_RNO_0_1_LC_15_3_1  (
            .in0(_gnd_net_),
            .in1(N__27221),
            .in2(N__27195),
            .in3(N__24939),
            .lcout(\QuadInstance4.Quad_RNO_0_3_1 ),
            .ltout(),
            .carryin(\QuadInstance4.un1_Quad_cry_0 ),
            .carryout(\QuadInstance4.un1_Quad_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_RNO_0_2_LC_15_3_2 .C_ON=1'b1;
    defparam \QuadInstance4.Quad_RNO_0_2_LC_15_3_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNO_0_2_LC_15_3_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance4.Quad_RNO_0_2_LC_15_3_2  (
            .in0(_gnd_net_),
            .in1(N__27178),
            .in2(N__27231),
            .in3(N__24936),
            .lcout(\QuadInstance4.Quad_RNO_0_4_2 ),
            .ltout(),
            .carryin(\QuadInstance4.un1_Quad_cry_1 ),
            .carryout(\QuadInstance4.un1_Quad_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_RNO_0_3_LC_15_3_3 .C_ON=1'b1;
    defparam \QuadInstance4.Quad_RNO_0_3_LC_15_3_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNO_0_3_LC_15_3_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance4.Quad_RNO_0_3_LC_15_3_3  (
            .in0(_gnd_net_),
            .in1(N__28043),
            .in2(N__27159),
            .in3(N__24933),
            .lcout(\QuadInstance4.Quad_RNO_0_4_3 ),
            .ltout(),
            .carryin(\QuadInstance4.un1_Quad_cry_2 ),
            .carryout(\QuadInstance4.un1_Quad_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_RNO_0_4_LC_15_3_4 .C_ON=1'b1;
    defparam \QuadInstance4.Quad_RNO_0_4_LC_15_3_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNO_0_4_LC_15_3_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance4.Quad_RNO_0_4_LC_15_3_4  (
            .in0(_gnd_net_),
            .in1(N__27528),
            .in2(N__27498),
            .in3(N__24918),
            .lcout(\QuadInstance4.Quad_RNO_0_4_4 ),
            .ltout(),
            .carryin(\QuadInstance4.un1_Quad_cry_3 ),
            .carryout(\QuadInstance4.un1_Quad_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_RNO_0_5_LC_15_3_5 .C_ON=1'b1;
    defparam \QuadInstance4.Quad_RNO_0_5_LC_15_3_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNO_0_5_LC_15_3_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance4.Quad_RNO_0_5_LC_15_3_5  (
            .in0(_gnd_net_),
            .in1(N__27053),
            .in2(N__27036),
            .in3(N__25062),
            .lcout(\QuadInstance4.Quad_RNO_0_4_5 ),
            .ltout(),
            .carryin(\QuadInstance4.un1_Quad_cry_4 ),
            .carryout(\QuadInstance4.un1_Quad_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_RNO_0_6_LC_15_3_6 .C_ON=1'b1;
    defparam \QuadInstance4.Quad_RNO_0_6_LC_15_3_6 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNO_0_6_LC_15_3_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance4.Quad_RNO_0_6_LC_15_3_6  (
            .in0(_gnd_net_),
            .in1(N__25087),
            .in2(N__25158),
            .in3(N__25059),
            .lcout(\QuadInstance4.Quad_RNO_0_4_6 ),
            .ltout(),
            .carryin(\QuadInstance4.un1_Quad_cry_5 ),
            .carryout(\QuadInstance4.un1_Quad_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_RNO_0_7_LC_15_3_7 .C_ON=1'b1;
    defparam \QuadInstance4.Quad_RNO_0_7_LC_15_3_7 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNO_0_7_LC_15_3_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance4.Quad_RNO_0_7_LC_15_3_7  (
            .in0(_gnd_net_),
            .in1(N__27648),
            .in2(N__25239),
            .in3(N__25056),
            .lcout(\QuadInstance4.Quad_RNO_0_4_7 ),
            .ltout(),
            .carryin(\QuadInstance4.un1_Quad_cry_6 ),
            .carryout(\QuadInstance4.un1_Quad_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_RNO_0_8_LC_15_4_0 .C_ON=1'b1;
    defparam \QuadInstance4.Quad_RNO_0_8_LC_15_4_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNO_0_8_LC_15_4_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance4.Quad_RNO_0_8_LC_15_4_0  (
            .in0(_gnd_net_),
            .in1(N__27264),
            .in2(N__27285),
            .in3(N__25053),
            .lcout(\QuadInstance4.Quad_RNO_0_4_8 ),
            .ltout(),
            .carryin(bfn_15_4_0_),
            .carryout(\QuadInstance4.un1_Quad_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_RNO_0_9_LC_15_4_1 .C_ON=1'b1;
    defparam \QuadInstance4.Quad_RNO_0_9_LC_15_4_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNO_0_9_LC_15_4_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance4.Quad_RNO_0_9_LC_15_4_1  (
            .in0(_gnd_net_),
            .in1(N__25348),
            .in2(N__25251),
            .in3(N__25035),
            .lcout(\QuadInstance4.Quad_RNO_0_4_9 ),
            .ltout(),
            .carryin(\QuadInstance4.un1_Quad_cry_8 ),
            .carryout(\QuadInstance4.un1_Quad_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_RNO_0_10_LC_15_4_2 .C_ON=1'b1;
    defparam \QuadInstance4.Quad_RNO_0_10_LC_15_4_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNO_0_10_LC_15_4_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance4.Quad_RNO_0_10_LC_15_4_2  (
            .in0(_gnd_net_),
            .in1(N__32867),
            .in2(N__25146),
            .in3(N__25032),
            .lcout(\QuadInstance4.Quad_RNO_0_4_10 ),
            .ltout(),
            .carryin(\QuadInstance4.un1_Quad_cry_9 ),
            .carryout(\QuadInstance4.un1_Quad_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_RNO_0_11_LC_15_4_3 .C_ON=1'b1;
    defparam \QuadInstance4.Quad_RNO_0_11_LC_15_4_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNO_0_11_LC_15_4_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance4.Quad_RNO_0_11_LC_15_4_3  (
            .in0(_gnd_net_),
            .in1(N__25108),
            .in2(N__25137),
            .in3(N__25029),
            .lcout(\QuadInstance4.Quad_RNO_0_4_11 ),
            .ltout(),
            .carryin(\QuadInstance4.un1_Quad_cry_10 ),
            .carryout(\QuadInstance4.un1_Quad_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_RNO_0_12_LC_15_4_4 .C_ON=1'b1;
    defparam \QuadInstance4.Quad_RNO_0_12_LC_15_4_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNO_0_12_LC_15_4_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance4.Quad_RNO_0_12_LC_15_4_4  (
            .in0(_gnd_net_),
            .in1(N__27027),
            .in2(N__27603),
            .in3(N__25026),
            .lcout(\QuadInstance4.Quad_RNO_0_4_12 ),
            .ltout(),
            .carryin(\QuadInstance4.un1_Quad_cry_11 ),
            .carryout(\QuadInstance4.un1_Quad_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_RNO_0_13_LC_15_4_5 .C_ON=1'b1;
    defparam \QuadInstance4.Quad_RNO_0_13_LC_15_4_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNO_0_13_LC_15_4_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance4.Quad_RNO_0_13_LC_15_4_5  (
            .in0(_gnd_net_),
            .in1(N__27569),
            .in2(N__27150),
            .in3(N__25023),
            .lcout(\QuadInstance4.Quad_RNO_0_4_13 ),
            .ltout(),
            .carryin(\QuadInstance4.un1_Quad_cry_12 ),
            .carryout(\QuadInstance4.un1_Quad_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_RNO_0_14_LC_15_4_6 .C_ON=1'b1;
    defparam \QuadInstance4.Quad_RNO_0_14_LC_15_4_6 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNO_0_14_LC_15_4_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance4.Quad_RNO_0_14_LC_15_4_6  (
            .in0(_gnd_net_),
            .in1(N__27141),
            .in2(N__29969),
            .in3(N__25188),
            .lcout(\QuadInstance4.Quad_RNO_0_4_14 ),
            .ltout(),
            .carryin(\QuadInstance4.un1_Quad_cry_13 ),
            .carryout(\QuadInstance4.un1_Quad_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_15_LC_15_4_7 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_15_LC_15_4_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance4.Quad_15_LC_15_4_7 .LUT_INIT=16'b1101000111100010;
    LogicCell40 \QuadInstance4.Quad_15_LC_15_4_7  (
            .in0(N__25185),
            .in1(N__29628),
            .in2(N__31916),
            .in3(N__25170),
            .lcout(dataRead4_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38705),
            .ce(),
            .sr(N__35716));
    defparam \QuadInstance0.Quad_6_LC_15_5_1 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_6_LC_15_5_1 .SEQ_MODE=4'b1000;
    defparam \QuadInstance0.Quad_6_LC_15_5_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance0.Quad_6_LC_15_5_1  (
            .in0(N__31107),
            .in1(N__33120),
            .in2(_gnd_net_),
            .in3(N__30243),
            .lcout(dataRead0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38697),
            .ce(),
            .sr(N__35723));
    defparam \QuadInstance4.Quad_6_LC_15_5_2 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_6_LC_15_5_2 .SEQ_MODE=4'b1000;
    defparam \QuadInstance4.Quad_6_LC_15_5_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance4.Quad_6_LC_15_5_2  (
            .in0(N__31108),
            .in1(N__29604),
            .in2(_gnd_net_),
            .in3(N__25167),
            .lcout(dataRead4_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38697),
            .ce(),
            .sr(N__35723));
    defparam \QuadInstance4.Quad_RNIL00S1_6_LC_15_5_3 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_RNIL00S1_6_LC_15_5_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNIL00S1_6_LC_15_5_3 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \QuadInstance4.Quad_RNIL00S1_6_LC_15_5_3  (
            .in0(N__29600),
            .in1(N__27423),
            .in2(N__25089),
            .in3(N__27342),
            .lcout(\QuadInstance4.Quad_RNIL00S1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_RNI06TL1_10_LC_15_5_4 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_RNI06TL1_10_LC_15_5_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNI06TL1_10_LC_15_5_4 .LUT_INIT=16'b1111000001010000;
    LogicCell40 \QuadInstance4.Quad_RNI06TL1_10_LC_15_5_4  (
            .in0(N__27343),
            .in1(N__32871),
            .in2(N__27444),
            .in3(N__29601),
            .lcout(\QuadInstance4.Quad_RNI06TL1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_RNI17TL1_11_LC_15_5_5 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_RNI17TL1_11_LC_15_5_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNI17TL1_11_LC_15_5_5 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \QuadInstance4.Quad_RNI17TL1_11_LC_15_5_5  (
            .in0(N__29602),
            .in1(N__27344),
            .in2(N__25115),
            .in3(N__27427),
            .lcout(\QuadInstance4.Quad_RNI17TL1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_11_LC_15_5_7 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_11_LC_15_5_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance4.Quad_11_LC_15_5_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance4.Quad_11_LC_15_5_7  (
            .in0(N__29603),
            .in1(N__36012),
            .in2(_gnd_net_),
            .in3(N__25128),
            .lcout(dataRead4_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38697),
            .ce(),
            .sr(N__35723));
    defparam OutReg_esr_RNO_4_6_LC_15_6_0.C_ON=1'b0;
    defparam OutReg_esr_RNO_4_6_LC_15_6_0.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_4_6_LC_15_6_0.LUT_INIT=16'b0011001100011101;
    LogicCell40 OutReg_esr_RNO_4_6_LC_15_6_0 (
            .in0(N__33970),
            .in1(N__28127),
            .in2(N__25088),
            .in3(N__27976),
            .lcout(),
            .ltout(OutReg_0_5_i_m3_ns_1_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_esr_RNO_2_6_LC_15_6_1.C_ON=1'b0;
    defparam OutReg_esr_RNO_2_6_LC_15_6_1.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_2_6_LC_15_6_1.LUT_INIT=16'b1010110000001111;
    LogicCell40 OutReg_esr_RNO_2_6_LC_15_6_1 (
            .in0(N__25310),
            .in1(N__25280),
            .in2(N__25254),
            .in3(N__38094),
            .lcout(OutReg_esr_RNO_2Z0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam quadWrite_4_LC_15_6_2.C_ON=1'b0;
    defparam quadWrite_4_LC_15_6_2.SEQ_MODE=4'b1000;
    defparam quadWrite_4_LC_15_6_2.LUT_INIT=16'b0010000000000000;
    LogicCell40 quadWrite_4_LC_15_6_2 (
            .in0(N__33856),
            .in1(N__33658),
            .in2(N__33447),
            .in3(N__33234),
            .lcout(quadWriteZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38691),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_RNIO30S1_9_LC_15_6_3 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_RNIO30S1_9_LC_15_6_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNIO30S1_9_LC_15_6_3 .LUT_INIT=16'b1010111100000000;
    LogicCell40 \QuadInstance4.Quad_RNIO30S1_9_LC_15_6_3  (
            .in0(N__29599),
            .in1(N__25349),
            .in2(N__27353),
            .in3(N__27439),
            .lcout(\QuadInstance4.Quad_RNIO30S1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwmWrite_fast_4_LC_15_6_4.C_ON=1'b0;
    defparam pwmWrite_fast_4_LC_15_6_4.SEQ_MODE=4'b1000;
    defparam pwmWrite_fast_4_LC_15_6_4.LUT_INIT=16'b0000001000000000;
    LogicCell40 pwmWrite_fast_4_LC_15_6_4 (
            .in0(N__33855),
            .in1(N__33657),
            .in2(N__33446),
            .in3(N__33233),
            .lcout(pwmWrite_fastZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38691),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_RNIM10S1_7_LC_15_6_6 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_RNIM10S1_7_LC_15_6_6 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNIM10S1_7_LC_15_6_6 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance4.Quad_RNIM10S1_7_LC_15_6_6  (
            .in0(N__27644),
            .in1(N__29598),
            .in2(N__27451),
            .in3(N__27338),
            .lcout(\QuadInstance4.Quad_RNIM10S1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_4_15_LC_15_7_0.C_ON=1'b0;
    defparam OutReg_ess_RNO_4_15_LC_15_7_0.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_4_15_LC_15_7_0.LUT_INIT=16'b0001110000011111;
    LogicCell40 OutReg_ess_RNO_4_15_LC_15_7_0 (
            .in0(N__25214),
            .in1(N__32908),
            .in2(N__32818),
            .in3(N__30581),
            .lcout(OutReg_0_5_i_m3_ns_1_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_RNO_0_15_LC_15_7_1 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_RNO_0_15_LC_15_7_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNO_0_15_LC_15_7_1 .LUT_INIT=16'b0110101001011010;
    LogicCell40 \QuadInstance0.Quad_RNO_0_15_LC_15_7_1  (
            .in0(N__30582),
            .in1(N__33111),
            .in2(N__34086),
            .in3(N__33944),
            .lcout(\QuadInstance0.un1_Quad_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_received_0_rep2_esr_LC_15_7_2.C_ON=1'b0;
    defparam data_received_0_rep2_esr_LC_15_7_2.SEQ_MODE=4'b1000;
    defparam data_received_0_rep2_esr_LC_15_7_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 data_received_0_rep2_esr_LC_15_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35086),
            .lcout(data_received_0_repZ0Z2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38683),
            .ce(N__26179),
            .sr(N__26157));
    defparam \QuadInstance0.Quad_RNIOMBH1_9_LC_15_7_3 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_RNIOMBH1_9_LC_15_7_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNIOMBH1_9_LC_15_7_3 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance0.Quad_RNIOMBH1_9_LC_15_7_3  (
            .in0(N__30161),
            .in1(N__33110),
            .in2(N__34085),
            .in3(N__33943),
            .lcout(\QuadInstance0.Quad_RNIOMBH1Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_received_0_rep1_esr_LC_15_7_4.C_ON=1'b0;
    defparam data_received_0_rep1_esr_LC_15_7_4.SEQ_MODE=4'b1000;
    defparam data_received_0_rep1_esr_LC_15_7_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 data_received_0_rep1_esr_LC_15_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35085),
            .lcout(data_received_0_repZ0Z1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38683),
            .ce(N__26179),
            .sr(N__26157));
    defparam data_received_fast_esr_0_LC_15_7_5.C_ON=1'b0;
    defparam data_received_fast_esr_0_LC_15_7_5.SEQ_MODE=4'b1000;
    defparam data_received_fast_esr_0_LC_15_7_5.LUT_INIT=16'b1010101010101010;
    LogicCell40 data_received_fast_esr_0_LC_15_7_5 (
            .in0(N__35088),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(data_received_fastZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38683),
            .ce(N__26179),
            .sr(N__26157));
    defparam data_received_esr_0_LC_15_7_6.C_ON=1'b0;
    defparam data_received_esr_0_LC_15_7_6.SEQ_MODE=4'b1000;
    defparam data_received_esr_0_LC_15_7_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 data_received_esr_0_LC_15_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35087),
            .lcout(data_receivedZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38683),
            .ce(N__26179),
            .sr(N__26157));
    defparam data_received_esr_1_LC_15_7_7.C_ON=1'b0;
    defparam data_received_esr_1_LC_15_7_7.SEQ_MODE=4'b1000;
    defparam data_received_esr_1_LC_15_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 data_received_esr_1_LC_15_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38100),
            .lcout(data_receivedZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38683),
            .ce(N__26179),
            .sr(N__26157));
    defparam OutReg_ess_RNO_2_9_LC_15_8_0.C_ON=1'b0;
    defparam OutReg_ess_RNO_2_9_LC_15_8_0.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_2_9_LC_15_8_0.LUT_INIT=16'b1000100011110011;
    LogicCell40 OutReg_ess_RNO_2_9_LC_15_8_0 (
            .in0(N__25544),
            .in1(N__38095),
            .in2(N__25518),
            .in3(N__25317),
            .lcout(),
            .ltout(OutReg_ess_RNO_2Z0Z_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_0_9_LC_15_8_1.C_ON=1'b0;
    defparam OutReg_ess_RNO_0_9_LC_15_8_1.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_0_9_LC_15_8_1.LUT_INIT=16'b1111110000110000;
    LogicCell40 OutReg_ess_RNO_0_9_LC_15_8_1 (
            .in0(_gnd_net_),
            .in1(N__37505),
            .in2(N__25485),
            .in3(N__25356),
            .lcout(OutReg_ess_RNO_0Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_3_9_LC_15_8_2.C_ON=1'b0;
    defparam OutReg_ess_RNO_3_9_LC_15_8_2.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_3_9_LC_15_8_2.LUT_INIT=16'b0101010100100111;
    LogicCell40 OutReg_ess_RNO_3_9_LC_15_8_2 (
            .in0(N__34742),
            .in1(N__25482),
            .in2(N__25452),
            .in3(N__34863),
            .lcout(),
            .ltout(OutReg_0_4_i_m3_ns_1_9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_1_9_LC_15_8_3.C_ON=1'b0;
    defparam OutReg_ess_RNO_1_9_LC_15_8_3.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_1_9_LC_15_8_3.LUT_INIT=16'b1010110000001111;
    LogicCell40 OutReg_ess_RNO_1_9_LC_15_8_3 (
            .in0(N__25414),
            .in1(N__25391),
            .in2(N__25359),
            .in3(N__37701),
            .lcout(OutReg_ess_RNO_1Z0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_4_9_LC_15_8_4.C_ON=1'b0;
    defparam OutReg_ess_RNO_4_9_LC_15_8_4.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_4_9_LC_15_8_4.LUT_INIT=16'b0101010100011011;
    LogicCell40 OutReg_ess_RNO_4_9_LC_15_8_4 (
            .in0(N__32810),
            .in1(N__30157),
            .in2(N__25350),
            .in3(N__32922),
            .lcout(OutReg_0_5_i_m3_ns_1_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_received_2_rep2_esr_LC_15_8_5.C_ON=1'b0;
    defparam data_received_2_rep2_esr_LC_15_8_5.SEQ_MODE=4'b1000;
    defparam data_received_2_rep2_esr_LC_15_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 data_received_2_rep2_esr_LC_15_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37507),
            .lcout(data_received_2_repZ0Z2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38675),
            .ce(N__26180),
            .sr(N__26155));
    defparam data_received_esr_2_LC_15_8_6.C_ON=1'b0;
    defparam data_received_esr_2_LC_15_8_6.SEQ_MODE=4'b1000;
    defparam data_received_esr_2_LC_15_8_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 data_received_esr_2_LC_15_8_6 (
            .in0(N__37506),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(data_receivedZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38675),
            .ce(N__26180),
            .sr(N__26155));
    defparam \QuadInstance4.Quad_13_LC_15_9_0 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_13_LC_15_9_0 .SEQ_MODE=4'b1000;
    defparam \QuadInstance4.Quad_13_LC_15_9_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance4.Quad_13_LC_15_9_0  (
            .in0(N__28703),
            .in1(N__29642),
            .in2(_gnd_net_),
            .in3(N__26130),
            .lcout(dataRead4_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38666),
            .ce(),
            .sr(N__35752));
    defparam \QuadInstance7.Quad_13_LC_15_9_1 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_13_LC_15_9_1 .SEQ_MODE=4'b1000;
    defparam \QuadInstance7.Quad_13_LC_15_9_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance7.Quad_13_LC_15_9_1  (
            .in0(N__28704),
            .in1(N__26040),
            .in2(_gnd_net_),
            .in3(N__26121),
            .lcout(dataRead7_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38666),
            .ce(),
            .sr(N__35752));
    defparam \QuadInstance4.Quad_3_LC_15_9_2 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_3_LC_15_9_2 .SEQ_MODE=4'b1000;
    defparam \QuadInstance4.Quad_3_LC_15_9_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance4.Quad_3_LC_15_9_2  (
            .in0(N__32020),
            .in1(N__29643),
            .in2(_gnd_net_),
            .in3(N__26079),
            .lcout(dataRead4_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38666),
            .ce(),
            .sr(N__35752));
    defparam \QuadInstance7.Quad_3_LC_15_9_3 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_3_LC_15_9_3 .SEQ_MODE=4'b1000;
    defparam \QuadInstance7.Quad_3_LC_15_9_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance7.Quad_3_LC_15_9_3  (
            .in0(N__32022),
            .in1(N__26041),
            .in2(_gnd_net_),
            .in3(N__26070),
            .lcout(dataRead7_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38666),
            .ce(),
            .sr(N__35752));
    defparam \QuadInstance7.Quad_1_LC_15_9_4 .C_ON=1'b0;
    defparam \QuadInstance7.Quad_1_LC_15_9_4 .SEQ_MODE=4'b1000;
    defparam \QuadInstance7.Quad_1_LC_15_9_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance7.Quad_1_LC_15_9_4  (
            .in0(N__26039),
            .in1(N__31256),
            .in2(_gnd_net_),
            .in3(N__25857),
            .lcout(dataRead7_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38666),
            .ce(),
            .sr(N__35752));
    defparam \QuadInstance5.Quad_3_LC_15_9_5 .C_ON=1'b0;
    defparam \QuadInstance5.Quad_3_LC_15_9_5 .SEQ_MODE=4'b1000;
    defparam \QuadInstance5.Quad_3_LC_15_9_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance5.Quad_3_LC_15_9_5  (
            .in0(N__32021),
            .in1(N__25801),
            .in2(_gnd_net_),
            .in3(N__25641),
            .lcout(dataRead5_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38666),
            .ce(),
            .sr(N__35752));
    defparam GB_BUFFER_RST_c_i_g_THRU_LUT4_0_LC_15_9_6.C_ON=1'b0;
    defparam GB_BUFFER_RST_c_i_g_THRU_LUT4_0_LC_15_9_6.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_RST_c_i_g_THRU_LUT4_0_LC_15_9_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_RST_c_i_g_THRU_LUT4_0_LC_15_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35828),
            .lcout(GB_BUFFER_RST_c_i_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_2_7_LC_15_10_0.C_ON=1'b0;
    defparam OutReg_ess_RNO_2_7_LC_15_10_0.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_2_7_LC_15_10_0.LUT_INIT=16'b1010000011011101;
    LogicCell40 OutReg_ess_RNO_2_7_LC_15_10_0 (
            .in0(N__38139),
            .in1(N__25608),
            .in2(N__25575),
            .in3(N__27669),
            .lcout(),
            .ltout(OutReg_ess_RNO_2Z0Z_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_0_7_LC_15_10_1.C_ON=1'b0;
    defparam OutReg_ess_RNO_0_7_LC_15_10_1.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_0_7_LC_15_10_1.LUT_INIT=16'b1111101001010000;
    LogicCell40 OutReg_ess_RNO_0_7_LC_15_10_1 (
            .in0(N__37537),
            .in1(_gnd_net_),
            .in2(N__26382),
            .in3(N__26235),
            .lcout(),
            .ltout(OutReg_ess_RNO_0Z0Z_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_7_LC_15_10_2.C_ON=1'b0;
    defparam OutReg_ess_7_LC_15_10_2.SEQ_MODE=4'b1001;
    defparam OutReg_ess_7_LC_15_10_2.LUT_INIT=16'b1010101010111000;
    LogicCell40 OutReg_ess_7_LC_15_10_2 (
            .in0(N__28314),
            .in1(N__38879),
            .in2(N__26379),
            .in3(N__37378),
            .lcout(OutRegZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38654),
            .ce(N__37241),
            .sr(N__37129));
    defparam OutReg_ess_RNO_3_7_LC_15_10_3.C_ON=1'b0;
    defparam OutReg_ess_RNO_3_7_LC_15_10_3.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_3_7_LC_15_10_3.LUT_INIT=16'b0000001111011101;
    LogicCell40 OutReg_ess_RNO_3_7_LC_15_10_3 (
            .in0(N__26376),
            .in1(N__34883),
            .in2(N__26340),
            .in3(N__34762),
            .lcout(),
            .ltout(OutReg_0_4_i_m3_ns_1_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_1_7_LC_15_10_4.C_ON=1'b0;
    defparam OutReg_ess_RNO_1_7_LC_15_10_4.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_1_7_LC_15_10_4.LUT_INIT=16'b1010110000001111;
    LogicCell40 OutReg_ess_RNO_1_7_LC_15_10_4 (
            .in0(N__26304),
            .in1(N__26270),
            .in2(N__26238),
            .in3(N__37744),
            .lcout(OutReg_ess_RNO_1Z0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_9_LC_15_10_5.C_ON=1'b0;
    defparam OutReg_ess_9_LC_15_10_5.SEQ_MODE=4'b1001;
    defparam OutReg_ess_9_LC_15_10_5.LUT_INIT=16'b1100110111001000;
    LogicCell40 OutReg_ess_9_LC_15_10_5 (
            .in0(N__37379),
            .in1(N__37263),
            .in2(N__38910),
            .in3(N__26229),
            .lcout(OutRegZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38654),
            .ce(N__37241),
            .sr(N__37129));
    defparam OutReg_esr_14_LC_15_11_0.C_ON=1'b0;
    defparam OutReg_esr_14_LC_15_11_0.SEQ_MODE=4'b1000;
    defparam OutReg_esr_14_LC_15_11_0.LUT_INIT=16'b1111000111100000;
    LogicCell40 OutReg_esr_14_LC_15_11_0 (
            .in0(N__38937),
            .in1(N__37380),
            .in2(N__26220),
            .in3(N__28146),
            .lcout(OutRegZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38644),
            .ce(N__37246),
            .sr(N__37132));
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_15_12_0 .C_ON=1'b0;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_15_12_0 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance3.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_15_12_0  (
            .in0(N__26190),
            .in1(N__26401),
            .in2(N__28437),
            .in3(N__26451),
            .lcout(\PWMInstance3.un1_PWMPulseWidthCount_0_I_15_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance3.periodCounter_RNI1D3C_2_LC_15_12_1 .C_ON=1'b0;
    defparam \PWMInstance3.periodCounter_RNI1D3C_2_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance3.periodCounter_RNI1D3C_2_LC_15_12_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \PWMInstance3.periodCounter_RNI1D3C_2_LC_15_12_1  (
            .in0(_gnd_net_),
            .in1(N__29154),
            .in2(_gnd_net_),
            .in3(N__28348),
            .lcout(),
            .ltout(\PWMInstance3.un1_periodCounter12_1_0_a2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance3.periodCounter_RNI83NV_4_LC_15_12_2 .C_ON=1'b0;
    defparam \PWMInstance3.periodCounter_RNI83NV_4_LC_15_12_2 .SEQ_MODE=4'b0000;
    defparam \PWMInstance3.periodCounter_RNI83NV_4_LC_15_12_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \PWMInstance3.periodCounter_RNI83NV_4_LC_15_12_2  (
            .in0(N__26493),
            .in1(N__29109),
            .in2(N__26460),
            .in3(N__26402),
            .lcout(\PWMInstance3.un1_periodCounter12_1_0_a2_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance3.PWMPulseWidthCount_esr_4_LC_15_12_3 .C_ON=1'b0;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_4_LC_15_12_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_4_LC_15_12_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \PWMInstance3.PWMPulseWidthCount_esr_4_LC_15_12_3  (
            .in0(N__36438),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PWMInstance3.PWMPulseWidthCountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38635),
            .ce(N__29298),
            .sr(N__35772));
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_15_12_5 .C_ON=1'b0;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_15_12_5 .SEQ_MODE=4'b0000;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_15_12_5 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance3.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_15_12_5  (
            .in0(N__26445),
            .in1(N__26492),
            .in2(N__28416),
            .in3(N__26439),
            .lcout(\PWMInstance3.un1_PWMPulseWidthCount_0_I_33_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance3.periodCounter_0_LC_15_13_0 .C_ON=1'b1;
    defparam \PWMInstance3.periodCounter_0_LC_15_13_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.periodCounter_0_LC_15_13_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance3.periodCounter_0_LC_15_13_0  (
            .in0(_gnd_net_),
            .in1(N__29055),
            .in2(N__26433),
            .in3(N__26432),
            .lcout(\PWMInstance3.periodCounterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_15_13_0_),
            .carryout(\PWMInstance3.un1_periodCounter_2_cry_0 ),
            .clk(N__38622),
            .ce(),
            .sr(N__35305));
    defparam \PWMInstance3.periodCounter_1_LC_15_13_1 .C_ON=1'b1;
    defparam \PWMInstance3.periodCounter_1_LC_15_13_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.periodCounter_1_LC_15_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance3.periodCounter_1_LC_15_13_1  (
            .in0(_gnd_net_),
            .in1(N__29039),
            .in2(_gnd_net_),
            .in3(N__26412),
            .lcout(\PWMInstance3.periodCounterZ0Z_1 ),
            .ltout(),
            .carryin(\PWMInstance3.un1_periodCounter_2_cry_0 ),
            .carryout(\PWMInstance3.un1_periodCounter_2_cry_1 ),
            .clk(N__38622),
            .ce(),
            .sr(N__35305));
    defparam \PWMInstance3.periodCounter_2_LC_15_13_2 .C_ON=1'b1;
    defparam \PWMInstance3.periodCounter_2_LC_15_13_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.periodCounter_2_LC_15_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance3.periodCounter_2_LC_15_13_2  (
            .in0(_gnd_net_),
            .in1(N__28350),
            .in2(_gnd_net_),
            .in3(N__26409),
            .lcout(\PWMInstance3.periodCounterZ0Z_2 ),
            .ltout(),
            .carryin(\PWMInstance3.un1_periodCounter_2_cry_1 ),
            .carryout(\PWMInstance3.un1_periodCounter_2_cry_2 ),
            .clk(N__38622),
            .ce(),
            .sr(N__35305));
    defparam \PWMInstance3.periodCounter_3_LC_15_13_3 .C_ON=1'b1;
    defparam \PWMInstance3.periodCounter_3_LC_15_13_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.periodCounter_3_LC_15_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance3.periodCounter_3_LC_15_13_3  (
            .in0(_gnd_net_),
            .in1(N__28367),
            .in2(_gnd_net_),
            .in3(N__26406),
            .lcout(\PWMInstance3.periodCounterZ0Z_3 ),
            .ltout(),
            .carryin(\PWMInstance3.un1_periodCounter_2_cry_2 ),
            .carryout(\PWMInstance3.un1_periodCounter_2_cry_3 ),
            .clk(N__38622),
            .ce(),
            .sr(N__35305));
    defparam \PWMInstance3.periodCounter_4_LC_15_13_4 .C_ON=1'b1;
    defparam \PWMInstance3.periodCounter_4_LC_15_13_4 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.periodCounter_4_LC_15_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance3.periodCounter_4_LC_15_13_4  (
            .in0(_gnd_net_),
            .in1(N__26403),
            .in2(_gnd_net_),
            .in3(N__26388),
            .lcout(\PWMInstance3.periodCounterZ0Z_4 ),
            .ltout(),
            .carryin(\PWMInstance3.un1_periodCounter_2_cry_3 ),
            .carryout(\PWMInstance3.un1_periodCounter_2_cry_4 ),
            .clk(N__38622),
            .ce(),
            .sr(N__35305));
    defparam \PWMInstance3.periodCounter_5_LC_15_13_5 .C_ON=1'b1;
    defparam \PWMInstance3.periodCounter_5_LC_15_13_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.periodCounter_5_LC_15_13_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance3.periodCounter_5_LC_15_13_5  (
            .in0(_gnd_net_),
            .in1(N__28436),
            .in2(_gnd_net_),
            .in3(N__26385),
            .lcout(\PWMInstance3.periodCounterZ0Z_5 ),
            .ltout(),
            .carryin(\PWMInstance3.un1_periodCounter_2_cry_4 ),
            .carryout(\PWMInstance3.un1_periodCounter_2_cry_5 ),
            .clk(N__38622),
            .ce(),
            .sr(N__35305));
    defparam \PWMInstance3.periodCounter_6_LC_15_13_6 .C_ON=1'b1;
    defparam \PWMInstance3.periodCounter_6_LC_15_13_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.periodCounter_6_LC_15_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance3.periodCounter_6_LC_15_13_6  (
            .in0(_gnd_net_),
            .in1(N__29481),
            .in2(_gnd_net_),
            .in3(N__26505),
            .lcout(\PWMInstance3.periodCounterZ0Z_6 ),
            .ltout(),
            .carryin(\PWMInstance3.un1_periodCounter_2_cry_5 ),
            .carryout(\PWMInstance3.un1_periodCounter_2_cry_6 ),
            .clk(N__38622),
            .ce(),
            .sr(N__35305));
    defparam \PWMInstance3.periodCounter_7_LC_15_13_7 .C_ON=1'b1;
    defparam \PWMInstance3.periodCounter_7_LC_15_13_7 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.periodCounter_7_LC_15_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance3.periodCounter_7_LC_15_13_7  (
            .in0(N__29765),
            .in1(N__29501),
            .in2(_gnd_net_),
            .in3(N__26502),
            .lcout(\PWMInstance3.periodCounterZ0Z_7 ),
            .ltout(),
            .carryin(\PWMInstance3.un1_periodCounter_2_cry_6 ),
            .carryout(\PWMInstance3.un1_periodCounter_2_cry_7 ),
            .clk(N__38622),
            .ce(),
            .sr(N__35305));
    defparam \PWMInstance3.periodCounter_8_LC_15_14_0 .C_ON=1'b1;
    defparam \PWMInstance3.periodCounter_8_LC_15_14_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.periodCounter_8_LC_15_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance3.periodCounter_8_LC_15_14_0  (
            .in0(_gnd_net_),
            .in1(N__29261),
            .in2(_gnd_net_),
            .in3(N__26499),
            .lcout(\PWMInstance3.periodCounterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_15_14_0_),
            .carryout(\PWMInstance3.un1_periodCounter_2_cry_8 ),
            .clk(N__38613),
            .ce(),
            .sr(N__35302));
    defparam \PWMInstance3.periodCounter_9_LC_15_14_1 .C_ON=1'b1;
    defparam \PWMInstance3.periodCounter_9_LC_15_14_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.periodCounter_9_LC_15_14_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance3.periodCounter_9_LC_15_14_1  (
            .in0(_gnd_net_),
            .in1(N__29243),
            .in2(_gnd_net_),
            .in3(N__26496),
            .lcout(\PWMInstance3.periodCounterZ0Z_9 ),
            .ltout(),
            .carryin(\PWMInstance3.un1_periodCounter_2_cry_8 ),
            .carryout(\PWMInstance3.un1_periodCounter_2_cry_9 ),
            .clk(N__38613),
            .ce(),
            .sr(N__35302));
    defparam \PWMInstance3.periodCounter_10_LC_15_14_2 .C_ON=1'b1;
    defparam \PWMInstance3.periodCounter_10_LC_15_14_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.periodCounter_10_LC_15_14_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance3.periodCounter_10_LC_15_14_2  (
            .in0(_gnd_net_),
            .in1(N__26491),
            .in2(_gnd_net_),
            .in3(N__26475),
            .lcout(\PWMInstance3.periodCounterZ0Z_10 ),
            .ltout(),
            .carryin(\PWMInstance3.un1_periodCounter_2_cry_9 ),
            .carryout(\PWMInstance3.un1_periodCounter_2_cry_10 ),
            .clk(N__38613),
            .ce(),
            .sr(N__35302));
    defparam \PWMInstance3.periodCounter_11_LC_15_14_3 .C_ON=1'b1;
    defparam \PWMInstance3.periodCounter_11_LC_15_14_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.periodCounter_11_LC_15_14_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance3.periodCounter_11_LC_15_14_3  (
            .in0(N__29766),
            .in1(N__28411),
            .in2(_gnd_net_),
            .in3(N__26472),
            .lcout(\PWMInstance3.periodCounterZ0Z_11 ),
            .ltout(),
            .carryin(\PWMInstance3.un1_periodCounter_2_cry_10 ),
            .carryout(\PWMInstance3.un1_periodCounter_2_cry_11 ),
            .clk(N__38613),
            .ce(),
            .sr(N__35302));
    defparam \PWMInstance3.periodCounter_12_LC_15_14_4 .C_ON=1'b1;
    defparam \PWMInstance3.periodCounter_12_LC_15_14_4 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.periodCounter_12_LC_15_14_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance3.periodCounter_12_LC_15_14_4  (
            .in0(N__29764),
            .in1(N__29108),
            .in2(_gnd_net_),
            .in3(N__26469),
            .lcout(\PWMInstance3.periodCounterZ0Z_12 ),
            .ltout(),
            .carryin(\PWMInstance3.un1_periodCounter_2_cry_11 ),
            .carryout(\PWMInstance3.un1_periodCounter_2_cry_12 ),
            .clk(N__38613),
            .ce(),
            .sr(N__35302));
    defparam \PWMInstance3.periodCounter_13_LC_15_14_5 .C_ON=1'b1;
    defparam \PWMInstance3.periodCounter_13_LC_15_14_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.periodCounter_13_LC_15_14_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance3.periodCounter_13_LC_15_14_5  (
            .in0(N__29767),
            .in1(N__29087),
            .in2(_gnd_net_),
            .in3(N__26466),
            .lcout(\PWMInstance3.periodCounterZ0Z_13 ),
            .ltout(),
            .carryin(\PWMInstance3.un1_periodCounter_2_cry_12 ),
            .carryout(\PWMInstance3.un1_periodCounter_2_cry_13 ),
            .clk(N__38613),
            .ce(),
            .sr(N__35302));
    defparam \PWMInstance3.periodCounter_14_LC_15_14_6 .C_ON=1'b1;
    defparam \PWMInstance3.periodCounter_14_LC_15_14_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.periodCounter_14_LC_15_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance3.periodCounter_14_LC_15_14_6  (
            .in0(_gnd_net_),
            .in1(N__29153),
            .in2(_gnd_net_),
            .in3(N__26463),
            .lcout(\PWMInstance3.periodCounterZ0Z_14 ),
            .ltout(),
            .carryin(\PWMInstance3.un1_periodCounter_2_cry_13 ),
            .carryout(\PWMInstance3.un1_periodCounter_2_cry_14 ),
            .clk(N__38613),
            .ce(),
            .sr(N__35302));
    defparam \PWMInstance3.periodCounter_15_LC_15_14_7 .C_ON=1'b1;
    defparam \PWMInstance3.periodCounter_15_LC_15_14_7 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.periodCounter_15_LC_15_14_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance3.periodCounter_15_LC_15_14_7  (
            .in0(_gnd_net_),
            .in1(N__29174),
            .in2(_gnd_net_),
            .in3(N__26715),
            .lcout(\PWMInstance3.periodCounterZ0Z_15 ),
            .ltout(),
            .carryin(\PWMInstance3.un1_periodCounter_2_cry_14 ),
            .carryout(\PWMInstance3.un1_periodCounter_2_cry_15 ),
            .clk(N__38613),
            .ce(),
            .sr(N__35302));
    defparam \PWMInstance3.periodCounter_16_LC_15_15_0 .C_ON=1'b0;
    defparam \PWMInstance3.periodCounter_16_LC_15_15_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.periodCounter_16_LC_15_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance3.periodCounter_16_LC_15_15_0  (
            .in0(N__29771),
            .in1(N__26704),
            .in2(_gnd_net_),
            .in3(N__26712),
            .lcout(\PWMInstance3.periodCounterZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38601),
            .ce(),
            .sr(N__35300));
    defparam \PWMInstance4.periodCounter_RNIQOSE_0_LC_15_16_0 .C_ON=1'b0;
    defparam \PWMInstance4.periodCounter_RNIQOSE_0_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance4.periodCounter_RNIQOSE_0_LC_15_16_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \PWMInstance4.periodCounter_RNIQOSE_0_LC_15_16_0  (
            .in0(N__26618),
            .in1(N__26684),
            .in2(N__26568),
            .in3(N__26663),
            .lcout(\PWMInstance4.un1_periodCounter12_1_0_a2_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_15_16_1 .C_ON=1'b0;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_15_16_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_15_16_1 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \PWMInstance4.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_15_16_1  (
            .in0(N__26662),
            .in1(N__26625),
            .in2(N__26814),
            .in3(N__26649),
            .lcout(\PWMInstance4.un1_PWMPulseWidthCount_0_I_1_c_RNO_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance4.PWMPulseWidthCount_esr_1_LC_15_16_3 .C_ON=1'b0;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_1_LC_15_16_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_1_LC_15_16_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \PWMInstance4.PWMPulseWidthCount_esr_1_LC_15_16_3  (
            .in0(N__31281),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PWMInstance4.PWMPulseWidthCountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38594),
            .ce(N__26934),
            .sr(N__35789));
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_15_16_4 .C_ON=1'b0;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_15_16_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_15_16_4 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \PWMInstance4.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_15_16_4  (
            .in0(N__26617),
            .in1(N__26592),
            .in2(N__26586),
            .in3(N__26993),
            .lcout(\PWMInstance4.un1_PWMPulseWidthCount_0_I_27_c_RNO_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance4.PWMPulseWidthCount_esr_6_LC_15_16_5 .C_ON=1'b0;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_6_LC_15_16_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_6_LC_15_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance4.PWMPulseWidthCount_esr_6_LC_15_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31118),
            .lcout(\PWMInstance4.PWMPulseWidthCountZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38594),
            .ce(N__26934),
            .sr(N__35789));
    defparam \PWMInstance4.PWMPulseWidthCount_esr_7_LC_15_16_6 .C_ON=1'b0;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_7_LC_15_16_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_7_LC_15_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance4.PWMPulseWidthCount_esr_7_LC_15_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29418),
            .lcout(\PWMInstance4.PWMPulseWidthCountZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38594),
            .ce(N__26934),
            .sr(N__35789));
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_15_16_7 .C_ON=1'b0;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_15_16_7 .SEQ_MODE=4'b0000;
    defparam \PWMInstance4.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_15_16_7 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance4.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_15_16_7  (
            .in0(N__26577),
            .in1(N__26563),
            .in2(N__26549),
            .in3(N__26526),
            .lcout(\PWMInstance4.un1_PWMPulseWidthCount_0_I_45_c_RNO_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance4.out_RNO_0_LC_15_17_0 .C_ON=1'b0;
    defparam \PWMInstance4.out_RNO_0_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance4.out_RNO_0_LC_15_17_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \PWMInstance4.out_RNO_0_LC_15_17_0  (
            .in0(N__26869),
            .in1(N__26904),
            .in2(N__26889),
            .in3(N__27008),
            .lcout(\PWMInstance4.un1_periodCounter12_1_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance4.clkCount_0_LC_15_17_1 .C_ON=1'b0;
    defparam \PWMInstance4.clkCount_0_LC_15_17_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.clkCount_0_LC_15_17_1 .LUT_INIT=16'b1010101000010001;
    LogicCell40 \PWMInstance4.clkCount_0_LC_15_17_1  (
            .in0(N__26975),
            .in1(N__26887),
            .in2(_gnd_net_),
            .in3(N__26870),
            .lcout(\PWMInstance4.clkCountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38583),
            .ce(),
            .sr(N__35793));
    defparam \PWMInstance4.periodCounter_RNIAN5D_16_LC_15_17_2 .C_ON=1'b0;
    defparam \PWMInstance4.periodCounter_RNIAN5D_16_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \PWMInstance4.periodCounter_RNIAN5D_16_LC_15_17_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \PWMInstance4.periodCounter_RNIAN5D_16_LC_15_17_2  (
            .in0(_gnd_net_),
            .in1(N__27007),
            .in2(_gnd_net_),
            .in3(N__26992),
            .lcout(\PWMInstance4.un1_periodCounter12_1_0_a2_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance4.clkCount_1_LC_15_17_3 .C_ON=1'b0;
    defparam \PWMInstance4.clkCount_1_LC_15_17_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance4.clkCount_1_LC_15_17_3 .LUT_INIT=16'b1001100110001000;
    LogicCell40 \PWMInstance4.clkCount_1_LC_15_17_3  (
            .in0(N__26976),
            .in1(N__26888),
            .in2(_gnd_net_),
            .in3(N__26871),
            .lcout(\PWMInstance4.clkCountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38583),
            .ce(),
            .sr(N__35793));
    defparam \PWMInstance4.PWMPulseWidthCount_esr_ctle_15_LC_15_17_4 .C_ON=1'b0;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_ctle_15_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance4.PWMPulseWidthCount_esr_ctle_15_LC_15_17_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \PWMInstance4.PWMPulseWidthCount_esr_ctle_15_LC_15_17_4  (
            .in0(_gnd_net_),
            .in1(N__35832),
            .in2(_gnd_net_),
            .in3(N__26974),
            .lcout(\PWMInstance4.pwmWrite_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance4.clkCount_RNI5QJC_0_LC_15_17_5 .C_ON=1'b0;
    defparam \PWMInstance4.clkCount_RNI5QJC_0_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \PWMInstance4.clkCount_RNI5QJC_0_LC_15_17_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \PWMInstance4.clkCount_RNI5QJC_0_LC_15_17_5  (
            .in0(N__26903),
            .in1(N__26883),
            .in2(_gnd_net_),
            .in3(N__26868),
            .lcout(\PWMInstance4.periodCounter12 ),
            .ltout(\PWMInstance4.periodCounter12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance4.periodCounter_RNII1V61_1_LC_15_17_6 .C_ON=1'b0;
    defparam \PWMInstance4.periodCounter_RNII1V61_1_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \PWMInstance4.periodCounter_RNII1V61_1_LC_15_17_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \PWMInstance4.periodCounter_RNII1V61_1_LC_15_17_6  (
            .in0(N__26833),
            .in1(N__26812),
            .in2(N__26793),
            .in3(N__26790),
            .lcout(),
            .ltout(\PWMInstance4.un1_periodCounter12_1_0_a2_0_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance4.periodCounter_RNIKFDB3_0_LC_15_17_7 .C_ON=1'b0;
    defparam \PWMInstance4.periodCounter_RNIKFDB3_0_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \PWMInstance4.periodCounter_RNIKFDB3_0_LC_15_17_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \PWMInstance4.periodCounter_RNIKFDB3_0_LC_15_17_7  (
            .in0(N__26784),
            .in1(N__26775),
            .in2(N__26769),
            .in3(N__26766),
            .lcout(\PWMInstance4.out_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance6.delayedCh_B_0_LC_15_18_5 .C_ON=1'b0;
    defparam \QuadInstance6.delayedCh_B_0_LC_15_18_5 .SEQ_MODE=4'b1000;
    defparam \QuadInstance6.delayedCh_B_0_LC_15_18_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \QuadInstance6.delayedCh_B_0_LC_15_18_5  (
            .in0(N__27120),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\QuadInstance6.delayedCh_BZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38573),
            .ce(),
            .sr(_gnd_net_));
    defparam PWM4_obufLegalizeSB_DFF_LC_15_20_0.C_ON=1'b0;
    defparam PWM4_obufLegalizeSB_DFF_LC_15_20_0.SEQ_MODE=4'b1000;
    defparam PWM4_obufLegalizeSB_DFF_LC_15_20_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 PWM4_obufLegalizeSB_DFF_LC_15_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PWM4_obufLegalizeSB_DFFNet),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36925),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.delayedCh_B_0_LC_16_2_4 .C_ON=1'b0;
    defparam \QuadInstance1.delayedCh_B_0_LC_16_2_4 .SEQ_MODE=4'b1000;
    defparam \QuadInstance1.delayedCh_B_0_LC_16_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance1.delayedCh_B_0_LC_16_2_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27084),
            .lcout(\QuadInstance1.delayedCh_BZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38721),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_4_5_LC_16_3_0.C_ON=1'b0;
    defparam OutReg_ess_RNO_4_5_LC_16_3_0.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_4_5_LC_16_3_0.LUT_INIT=16'b0001110000011111;
    LogicCell40 OutReg_ess_RNO_4_5_LC_16_3_0 (
            .in0(N__27052),
            .in1(N__28008),
            .in2(N__28139),
            .in3(N__34114),
            .lcout(OutReg_0_5_i_m3_ns_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_5_LC_16_3_2 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_5_LC_16_3_2 .SEQ_MODE=4'b1000;
    defparam \QuadInstance4.Quad_5_LC_16_3_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance4.Quad_5_LC_16_3_2  (
            .in0(N__29633),
            .in1(N__36347),
            .in2(_gnd_net_),
            .in3(N__27060),
            .lcout(dataRead4_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38718),
            .ce(),
            .sr(N__35717));
    defparam \QuadInstance4.Quad_RNIKVVR1_5_LC_16_3_3 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_RNIKVVR1_5_LC_16_3_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNIKVVR1_5_LC_16_3_3 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance4.Quad_RNIKVVR1_5_LC_16_3_3  (
            .in0(N__27054),
            .in1(N__29629),
            .in2(N__27445),
            .in3(N__27351),
            .lcout(\QuadInstance4.Quad_RNIKVVR1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_RNI28TL1_12_LC_16_3_4 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_RNI28TL1_12_LC_16_3_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNI28TL1_12_LC_16_3_4 .LUT_INIT=16'b1100010011000100;
    LogicCell40 \QuadInstance4.Quad_RNI28TL1_12_LC_16_3_4  (
            .in0(N__27352),
            .in1(N__27431),
            .in2(N__29652),
            .in3(N__27599),
            .lcout(\QuadInstance4.Quad_RNI28TL1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_esr_RNO_4_2_LC_16_4_0.C_ON=1'b0;
    defparam OutReg_esr_RNO_4_2_LC_16_4_0.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_4_2_LC_16_4_0.LUT_INIT=16'b0011001100011101;
    LogicCell40 OutReg_esr_RNO_4_2_LC_16_4_0 (
            .in0(N__32650),
            .in1(N__28132),
            .in2(N__27180),
            .in3(N__27989),
            .lcout(OutReg_0_5_i_m3_ns_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_2_LC_16_4_1 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_2_LC_16_4_1 .SEQ_MODE=4'b1000;
    defparam \QuadInstance0.Quad_2_LC_16_4_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance0.Quad_2_LC_16_4_1  (
            .in0(N__31585),
            .in1(N__33130),
            .in2(_gnd_net_),
            .in3(N__29877),
            .lcout(dataRead0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38711),
            .ce(),
            .sr(N__35724));
    defparam \QuadInstance4.delayedCh_A_RNIS1AU_2_LC_16_4_2 .C_ON=1'b0;
    defparam \QuadInstance4.delayedCh_A_RNIS1AU_2_LC_16_4_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.delayedCh_A_RNIS1AU_2_LC_16_4_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \QuadInstance4.delayedCh_A_RNIS1AU_2_LC_16_4_2  (
            .in0(N__27459),
            .in1(N__27474),
            .in2(N__29907),
            .in3(N__27134),
            .lcout(\QuadInstance4.count_enable ),
            .ltout(\QuadInstance4.count_enable_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_RNIHSVR1_2_LC_16_4_3 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_RNIHSVR1_2_LC_16_4_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNIHSVR1_2_LC_16_4_3 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance4.Quad_RNIHSVR1_2_LC_16_4_3  (
            .in0(N__27179),
            .in1(N__29622),
            .in2(N__27234),
            .in3(N__27331),
            .lcout(\QuadInstance4.Quad_RNIHSVR1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_RNIGRVR1_1_LC_16_4_5 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_RNIGRVR1_1_LC_16_4_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNIGRVR1_1_LC_16_4_5 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance4.Quad_RNIGRVR1_1_LC_16_4_5  (
            .in0(N__27222),
            .in1(N__29621),
            .in2(N__27440),
            .in3(N__27330),
            .lcout(\QuadInstance4.Quad_RNIGRVR1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_2_LC_16_4_6 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_2_LC_16_4_6 .SEQ_MODE=4'b1000;
    defparam \QuadInstance4.Quad_2_LC_16_4_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance4.Quad_2_LC_16_4_6  (
            .in0(N__29624),
            .in1(N__31586),
            .in2(_gnd_net_),
            .in3(N__27186),
            .lcout(dataRead4_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38711),
            .ce(),
            .sr(N__35724));
    defparam \QuadInstance4.Quad_RNIITVR1_3_LC_16_4_7 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_RNIITVR1_3_LC_16_4_7 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNIITVR1_3_LC_16_4_7 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance4.Quad_RNIITVR1_3_LC_16_4_7  (
            .in0(N__28044),
            .in1(N__29623),
            .in2(N__27441),
            .in3(N__27332),
            .lcout(\QuadInstance4.Quad_RNIITVR1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.delayedCh_B_2_LC_16_5_0 .C_ON=1'b0;
    defparam \QuadInstance4.delayedCh_B_2_LC_16_5_0 .SEQ_MODE=4'b1000;
    defparam \QuadInstance4.delayedCh_B_2_LC_16_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance4.delayedCh_B_2_LC_16_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29906),
            .lcout(\QuadInstance4.delayedCh_BZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38706),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_RNI39TL1_13_LC_16_5_1 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_RNI39TL1_13_LC_16_5_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNI39TL1_13_LC_16_5_1 .LUT_INIT=16'b1010000011110000;
    LogicCell40 \QuadInstance4.Quad_RNI39TL1_13_LC_16_5_1  (
            .in0(N__29589),
            .in1(N__27570),
            .in2(N__27443),
            .in3(N__27346),
            .lcout(\QuadInstance4.Quad_RNI39TL1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_RNI4ATL1_14_LC_16_5_2 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_RNI4ATL1_14_LC_16_5_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNI4ATL1_14_LC_16_5_2 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \QuadInstance4.Quad_RNI4ATL1_14_LC_16_5_2  (
            .in0(N__27347),
            .in1(N__29590),
            .in2(N__29965),
            .in3(N__27422),
            .lcout(\QuadInstance4.Quad_RNI4ATL1Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.delayedCh_B_RNISS9M_2_LC_16_5_3 .C_ON=1'b0;
    defparam \QuadInstance4.delayedCh_B_RNISS9M_2_LC_16_5_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.delayedCh_B_RNISS9M_2_LC_16_5_3 .LUT_INIT=16'b0000110011000000;
    LogicCell40 \QuadInstance4.delayedCh_B_RNISS9M_2_LC_16_5_3  (
            .in0(_gnd_net_),
            .in1(N__34496),
            .in2(N__27135),
            .in3(N__27472),
            .lcout(\QuadInstance4.un1_count_enable_i_a2_0_1 ),
            .ltout(\QuadInstance4.un1_count_enable_i_a2_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_RNIJUVR1_4_LC_16_5_4 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_RNIJUVR1_4_LC_16_5_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNIJUVR1_4_LC_16_5_4 .LUT_INIT=16'b1100111100000000;
    LogicCell40 \QuadInstance4.Quad_RNIJUVR1_4_LC_16_5_4  (
            .in0(N__27527),
            .in1(N__29587),
            .in2(N__27501),
            .in3(N__27415),
            .lcout(\QuadInstance4.Quad_RNIJUVR1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.delayedCh_A_1_LC_16_5_5 .C_ON=1'b0;
    defparam \QuadInstance4.delayedCh_A_1_LC_16_5_5 .SEQ_MODE=4'b1000;
    defparam \QuadInstance4.delayedCh_A_1_LC_16_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance4.delayedCh_A_1_LC_16_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27486),
            .lcout(\QuadInstance4.delayedCh_AZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38706),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.delayedCh_A_2_LC_16_5_6 .C_ON=1'b0;
    defparam \QuadInstance4.delayedCh_A_2_LC_16_5_6 .SEQ_MODE=4'b1000;
    defparam \QuadInstance4.delayedCh_A_2_LC_16_5_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \QuadInstance4.delayedCh_A_2_LC_16_5_6  (
            .in0(N__27473),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\QuadInstance4.delayedCh_AZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38706),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.Quad_RNIN20S1_8_LC_16_5_7 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_RNIN20S1_8_LC_16_5_7 .SEQ_MODE=4'b0000;
    defparam \QuadInstance4.Quad_RNIN20S1_8_LC_16_5_7 .LUT_INIT=16'b1010000011110000;
    LogicCell40 \QuadInstance4.Quad_RNIN20S1_8_LC_16_5_7  (
            .in0(N__29588),
            .in1(N__27263),
            .in2(N__27442),
            .in3(N__27345),
            .lcout(\QuadInstance4.Quad_RNIN20S1Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_esr_RNO_4_8_LC_16_6_0.C_ON=1'b0;
    defparam OutReg_esr_RNO_4_8_LC_16_6_0.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_4_8_LC_16_6_0.LUT_INIT=16'b0011001100011101;
    LogicCell40 OutReg_esr_RNO_4_8_LC_16_6_0 (
            .in0(N__30193),
            .in1(N__32835),
            .in2(N__27259),
            .in3(N__32945),
            .lcout(OutReg_0_5_i_m3_ns_1_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_8_LC_16_6_1 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_8_LC_16_6_1 .SEQ_MODE=4'b1000;
    defparam \QuadInstance0.Quad_8_LC_16_6_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance0.Quad_8_LC_16_6_1  (
            .in0(N__33102),
            .in1(N__28990),
            .in2(_gnd_net_),
            .in3(N__30171),
            .lcout(dataRead0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38698),
            .ce(),
            .sr(N__35740));
    defparam \QuadInstance4.Quad_8_LC_16_6_2 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_8_LC_16_6_2 .SEQ_MODE=4'b1000;
    defparam \QuadInstance4.Quad_8_LC_16_6_2 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \QuadInstance4.Quad_8_LC_16_6_2  (
            .in0(N__28991),
            .in1(_gnd_net_),
            .in2(N__27276),
            .in3(N__29619),
            .lcout(dataRead4_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38698),
            .ce(),
            .sr(N__35740));
    defparam \QuadInstance0.Quad_RNINLBH1_8_LC_16_6_3 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_RNINLBH1_8_LC_16_6_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNINLBH1_8_LC_16_6_3 .LUT_INIT=16'b1010000011110000;
    LogicCell40 \QuadInstance0.Quad_RNINLBH1_8_LC_16_6_3  (
            .in0(N__33101),
            .in1(N__30194),
            .in2(N__34081),
            .in3(N__33942),
            .lcout(\QuadInstance0.Quad_RNINLBH1Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_RNIMKBH1_7_LC_16_6_4 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_RNIMKBH1_7_LC_16_6_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNIMKBH1_7_LC_16_6_4 .LUT_INIT=16'b1100111100000000;
    LogicCell40 \QuadInstance0.Quad_RNIMKBH1_7_LC_16_6_4  (
            .in0(N__30227),
            .in1(N__33100),
            .in2(N__33950),
            .in3(N__34061),
            .lcout(\QuadInstance0.Quad_RNIMKBH1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_4_7_LC_16_6_5.C_ON=1'b0;
    defparam OutReg_ess_RNO_4_7_LC_16_6_5.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_4_7_LC_16_6_5.LUT_INIT=16'b0001101000011111;
    LogicCell40 OutReg_ess_RNO_4_7_LC_16_6_5 (
            .in0(N__32946),
            .in1(N__27640),
            .in2(N__32841),
            .in3(N__30226),
            .lcout(OutReg_0_5_i_m3_ns_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_7_LC_16_6_6 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_7_LC_16_6_6 .SEQ_MODE=4'b1000;
    defparam \QuadInstance0.Quad_7_LC_16_6_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance0.Quad_7_LC_16_6_6  (
            .in0(N__29426),
            .in1(N__33103),
            .in2(_gnd_net_),
            .in3(N__30204),
            .lcout(dataRead0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38698),
            .ce(),
            .sr(N__35740));
    defparam \QuadInstance4.Quad_7_LC_16_6_7 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_7_LC_16_6_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance4.Quad_7_LC_16_6_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance4.Quad_7_LC_16_6_7  (
            .in0(N__29618),
            .in1(N__29427),
            .in2(_gnd_net_),
            .in3(N__27657),
            .lcout(dataRead4_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38698),
            .ce(),
            .sr(N__35740));
    defparam OutReg_esr_RNO_4_12_LC_16_7_0.C_ON=1'b0;
    defparam OutReg_esr_RNO_4_12_LC_16_7_0.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_4_12_LC_16_7_0.LUT_INIT=16'b0000010110111011;
    LogicCell40 OutReg_esr_RNO_4_12_LC_16_7_0 (
            .in0(N__32910),
            .in1(N__30049),
            .in2(N__27595),
            .in3(N__32801),
            .lcout(OutReg_0_5_i_m3_ns_1_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_12_LC_16_7_1 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_12_LC_16_7_1 .SEQ_MODE=4'b1000;
    defparam \QuadInstance0.Quad_12_LC_16_7_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance0.Quad_12_LC_16_7_1  (
            .in0(N__33115),
            .in1(N__28861),
            .in2(_gnd_net_),
            .in3(N__30024),
            .lcout(dataRead0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38692),
            .ce(),
            .sr(N__35748));
    defparam \QuadInstance4.Quad_12_LC_16_7_2 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_12_LC_16_7_2 .SEQ_MODE=4'b1000;
    defparam \QuadInstance4.Quad_12_LC_16_7_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance4.Quad_12_LC_16_7_2  (
            .in0(N__28862),
            .in1(N__29620),
            .in2(_gnd_net_),
            .in3(N__27612),
            .lcout(dataRead4_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38692),
            .ce(),
            .sr(N__35748));
    defparam \QuadInstance0.Quad_RNI2N8Q1_12_LC_16_7_3 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_RNI2N8Q1_12_LC_16_7_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNI2N8Q1_12_LC_16_7_3 .LUT_INIT=16'b1010000011110000;
    LogicCell40 \QuadInstance0.Quad_RNI2N8Q1_12_LC_16_7_3  (
            .in0(N__33113),
            .in1(N__30053),
            .in2(N__34087),
            .in3(N__33945),
            .lcout(\QuadInstance0.Quad_RNI2N8Q1Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_RNI1M8Q1_11_LC_16_7_4 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_RNI1M8Q1_11_LC_16_7_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNI1M8Q1_11_LC_16_7_4 .LUT_INIT=16'b1100111100000000;
    LogicCell40 \QuadInstance0.Quad_RNI1M8Q1_11_LC_16_7_4  (
            .in0(N__30099),
            .in1(N__33112),
            .in2(N__33951),
            .in3(N__34077),
            .lcout(\QuadInstance0.Quad_RNI1M8Q1Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_RNI3O8Q1_13_LC_16_7_5 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_RNI3O8Q1_13_LC_16_7_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNI3O8Q1_13_LC_16_7_5 .LUT_INIT=16'b1011000010110000;
    LogicCell40 \QuadInstance0.Quad_RNI3O8Q1_13_LC_16_7_5  (
            .in0(N__33114),
            .in1(N__33949),
            .in2(N__34088),
            .in3(N__30013),
            .lcout(\QuadInstance0.Quad_RNI3O8Q1Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_4_13_LC_16_7_6.C_ON=1'b0;
    defparam OutReg_ess_RNO_4_13_LC_16_7_6.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_4_13_LC_16_7_6.LUT_INIT=16'b0001000110101111;
    LogicCell40 OutReg_ess_RNO_4_13_LC_16_7_6 (
            .in0(N__32909),
            .in1(N__27565),
            .in2(N__30015),
            .in3(N__32800),
            .lcout(OutReg_0_5_i_m3_ns_1_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_13_LC_16_7_7 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_13_LC_16_7_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance0.Quad_13_LC_16_7_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \QuadInstance0.Quad_13_LC_16_7_7  (
            .in0(N__33116),
            .in1(N__28727),
            .in2(_gnd_net_),
            .in3(N__29988),
            .lcout(dataRead0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38692),
            .ce(),
            .sr(N__35748));
    defparam OutReg_ess_RNO_4_3_LC_16_8_0.C_ON=1'b0;
    defparam OutReg_ess_RNO_4_3_LC_16_8_0.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_4_3_LC_16_8_0.LUT_INIT=16'b0101010100011011;
    LogicCell40 OutReg_ess_RNO_4_3_LC_16_8_0 (
            .in0(N__28128),
            .in1(N__34217),
            .in2(N__28042),
            .in3(N__27977),
            .lcout(),
            .ltout(OutReg_0_5_i_m3_ns_1_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_2_3_LC_16_8_1.C_ON=1'b0;
    defparam OutReg_ess_RNO_2_3_LC_16_8_1.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_2_3_LC_16_8_1.LUT_INIT=16'b1100101000001111;
    LogicCell40 OutReg_ess_RNO_2_3_LC_16_8_1 (
            .in0(N__27913),
            .in1(N__27879),
            .in2(N__27846),
            .in3(N__38096),
            .lcout(OutReg_ess_RNO_2Z0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_1_3_LC_16_8_2.C_ON=1'b0;
    defparam OutReg_ess_RNO_1_3_LC_16_8_2.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_1_3_LC_16_8_2.LUT_INIT=16'b1100000010111011;
    LogicCell40 OutReg_ess_RNO_1_3_LC_16_8_2 (
            .in0(N__27843),
            .in1(N__37702),
            .in2(N__27816),
            .in3(N__27780),
            .lcout(),
            .ltout(OutReg_ess_RNO_1Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_0_3_LC_16_8_3.C_ON=1'b0;
    defparam OutReg_ess_RNO_0_3_LC_16_8_3.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_0_3_LC_16_8_3.LUT_INIT=16'b1111001111000000;
    LogicCell40 OutReg_ess_RNO_0_3_LC_16_8_3 (
            .in0(_gnd_net_),
            .in1(N__37511),
            .in2(N__27771),
            .in3(N__27768),
            .lcout(),
            .ltout(OutReg_ess_RNO_0Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_3_LC_16_8_4.C_ON=1'b0;
    defparam OutReg_ess_3_LC_16_8_4.SEQ_MODE=4'b1001;
    defparam OutReg_ess_3_LC_16_8_4.LUT_INIT=16'b1010101010111000;
    LogicCell40 OutReg_ess_3_LC_16_8_4 (
            .in0(N__30474),
            .in1(N__38947),
            .in2(N__27762),
            .in3(N__37385),
            .lcout(OutRegZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38684),
            .ce(N__37250),
            .sr(N__37136));
    defparam OutReg_ess_4_LC_16_8_5.C_ON=1'b0;
    defparam OutReg_ess_4_LC_16_8_5.SEQ_MODE=4'b1001;
    defparam OutReg_ess_4_LC_16_8_5.LUT_INIT=16'b1100110111001000;
    LogicCell40 OutReg_ess_4_LC_16_8_5 (
            .in0(N__37386),
            .in1(N__27759),
            .in2(N__38952),
            .in3(N__27753),
            .lcout(OutRegZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38684),
            .ce(N__37250),
            .sr(N__37136));
    defparam OutReg_esr_RNO_1_6_LC_16_9_0.C_ON=1'b0;
    defparam OutReg_esr_RNO_1_6_LC_16_9_0.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_1_6_LC_16_9_0.LUT_INIT=16'b1000100011110011;
    LogicCell40 OutReg_esr_RNO_1_6_LC_16_9_0 (
            .in0(N__27741),
            .in1(N__37703),
            .in2(N__27708),
            .in3(N__28233),
            .lcout(),
            .ltout(OutReg_esr_RNO_1Z0Z_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_esr_RNO_0_6_LC_16_9_1.C_ON=1'b0;
    defparam OutReg_esr_RNO_0_6_LC_16_9_1.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_0_6_LC_16_9_1.LUT_INIT=16'b1111001111000000;
    LogicCell40 OutReg_esr_RNO_0_6_LC_16_9_1 (
            .in0(_gnd_net_),
            .in1(N__37521),
            .in2(N__28332),
            .in3(N__28329),
            .lcout(),
            .ltout(OutReg_esr_RNO_0Z0Z_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_esr_6_LC_16_9_2.C_ON=1'b0;
    defparam OutReg_esr_6_LC_16_9_2.SEQ_MODE=4'b1000;
    defparam OutReg_esr_6_LC_16_9_2.LUT_INIT=16'b1100110011011000;
    LogicCell40 OutReg_esr_6_LC_16_9_2 (
            .in0(N__38933),
            .in1(N__36666),
            .in2(N__28317),
            .in3(N__37351),
            .lcout(OutRegZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38676),
            .ce(N__37244),
            .sr(N__37131));
    defparam OutReg_esr_RNO_3_6_LC_16_9_3.C_ON=1'b0;
    defparam OutReg_esr_RNO_3_6_LC_16_9_3.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_3_6_LC_16_9_3.LUT_INIT=16'b0000001111011101;
    LogicCell40 OutReg_esr_RNO_3_6_LC_16_9_3 (
            .in0(N__28304),
            .in1(N__34895),
            .in2(N__28269),
            .in3(N__34761),
            .lcout(OutReg_0_4_i_m3_ns_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_received_esr_RNIA81U_3_LC_16_10_0.C_ON=1'b0;
    defparam data_received_esr_RNIA81U_3_LC_16_10_0.SEQ_MODE=4'b0000;
    defparam data_received_esr_RNIA81U_3_LC_16_10_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 data_received_esr_RNIA81U_3_LC_16_10_0 (
            .in0(N__30634),
            .in1(N__37512),
            .in2(N__38137),
            .in3(N__37704),
            .lcout(OutReg_0_sqmuxa_0_a2_3_a2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pwmWrite_2_LC_16_10_1.C_ON=1'b0;
    defparam pwmWrite_2_LC_16_10_1.SEQ_MODE=4'b1000;
    defparam pwmWrite_2_LC_16_10_1.LUT_INIT=16'b0000010000000000;
    LogicCell40 pwmWrite_2_LC_16_10_1 (
            .in0(N__33850),
            .in1(N__33660),
            .in2(N__33463),
            .in3(N__33214),
            .lcout(pwmWriteZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38667),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_esr_RNO_4_14_LC_16_10_3.C_ON=1'b0;
    defparam OutReg_esr_RNO_4_14_LC_16_10_3.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_4_14_LC_16_10_3.LUT_INIT=16'b0011001100011101;
    LogicCell40 OutReg_esr_RNO_4_14_LC_16_10_3 (
            .in0(N__34251),
            .in1(N__32830),
            .in2(N__29970),
            .in3(N__32947),
            .lcout(),
            .ltout(OutReg_0_5_i_m3_ns_1_14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_esr_RNO_2_14_LC_16_10_4.C_ON=1'b0;
    defparam OutReg_esr_RNO_2_14_LC_16_10_4.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_2_14_LC_16_10_4.LUT_INIT=16'b1100101000001111;
    LogicCell40 OutReg_esr_RNO_2_14_LC_16_10_4 (
            .in0(N__28227),
            .in1(N__28191),
            .in2(N__28161),
            .in3(N__38113),
            .lcout(),
            .ltout(OutReg_esr_RNO_2Z0Z_14_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_esr_RNO_0_14_LC_16_10_5.C_ON=1'b0;
    defparam OutReg_esr_RNO_0_14_LC_16_10_5.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_0_14_LC_16_10_5.LUT_INIT=16'b1111101001010000;
    LogicCell40 OutReg_esr_RNO_0_14_LC_16_10_5 (
            .in0(N__37513),
            .in1(_gnd_net_),
            .in2(N__28158),
            .in3(N__28155),
            .lcout(OutReg_esr_RNO_0Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.PWMPulseWidthCount_esr_12_LC_16_11_0 .C_ON=1'b0;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_12_LC_16_11_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_12_LC_16_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance2.PWMPulseWidthCount_esr_12_LC_16_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28819),
            .lcout(\PWMInstance2.PWMPulseWidthCountZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38655),
            .ce(N__35854),
            .sr(N__35773));
    defparam \PWMInstance2.PWMPulseWidthCount_esr_13_LC_16_11_1 .C_ON=1'b0;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_13_LC_16_11_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_13_LC_16_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance2.PWMPulseWidthCount_esr_13_LC_16_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28699),
            .lcout(\PWMInstance2.PWMPulseWidthCountZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38655),
            .ce(N__35854),
            .sr(N__35773));
    defparam \PWMInstance2.PWMPulseWidthCount_esr_8_LC_16_11_2 .C_ON=1'b0;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_8_LC_16_11_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_8_LC_16_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance2.PWMPulseWidthCount_esr_8_LC_16_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28972),
            .lcout(\PWMInstance2.PWMPulseWidthCountZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38655),
            .ce(N__35854),
            .sr(N__35773));
    defparam \PWMInstance2.PWMPulseWidthCount_esr_9_LC_16_11_3 .C_ON=1'b0;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_9_LC_16_11_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_9_LC_16_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance2.PWMPulseWidthCount_esr_9_LC_16_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28506),
            .lcout(\PWMInstance2.PWMPulseWidthCountZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38655),
            .ce(N__35854),
            .sr(N__35773));
    defparam \PWMInstance2.PWMPulseWidthCount_esr_7_LC_16_11_4 .C_ON=1'b0;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_7_LC_16_11_4 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_7_LC_16_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance2.PWMPulseWidthCount_esr_7_LC_16_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29392),
            .lcout(\PWMInstance2.PWMPulseWidthCountZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38655),
            .ce(N__35854),
            .sr(N__35773));
    defparam \PWMInstance3.PWMPulseWidthCount_esr_12_LC_16_12_0 .C_ON=1'b0;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_12_LC_16_12_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_12_LC_16_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance3.PWMPulseWidthCount_esr_12_LC_16_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28871),
            .lcout(\PWMInstance3.PWMPulseWidthCountZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38645),
            .ce(N__29319),
            .sr(N__35776));
    defparam \PWMInstance3.PWMPulseWidthCount_esr_13_LC_16_12_1 .C_ON=1'b0;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_13_LC_16_12_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_13_LC_16_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance3.PWMPulseWidthCount_esr_13_LC_16_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28724),
            .lcout(\PWMInstance3.PWMPulseWidthCountZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38645),
            .ce(N__29319),
            .sr(N__35776));
    defparam \PWMInstance3.PWMPulseWidthCount_esr_9_LC_16_12_3 .C_ON=1'b0;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_9_LC_16_12_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_9_LC_16_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance3.PWMPulseWidthCount_esr_9_LC_16_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28541),
            .lcout(\PWMInstance3.PWMPulseWidthCountZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38645),
            .ce(N__29319),
            .sr(N__35776));
    defparam \PWMInstance3.periodCounter_RNINK9L_3_LC_16_13_0 .C_ON=1'b0;
    defparam \PWMInstance3.periodCounter_RNINK9L_3_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance3.periodCounter_RNINK9L_3_LC_16_13_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \PWMInstance3.periodCounter_RNINK9L_3_LC_16_13_0  (
            .in0(N__29242),
            .in1(N__28435),
            .in2(N__28415),
            .in3(N__28366),
            .lcout(\PWMInstance3.un1_periodCounter12_1_0_a2_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_16_13_1 .C_ON=1'b0;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_16_13_1 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance3.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_16_13_1  (
            .in0(N__28380),
            .in1(N__29181),
            .in2(N__28368),
            .in3(N__28349),
            .lcout(\PWMInstance3.un1_PWMPulseWidthCount_0_I_9_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance3.PWMPulseWidthCount_esr_2_LC_16_13_2 .C_ON=1'b0;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_2_LC_16_13_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_2_LC_16_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance3.PWMPulseWidthCount_esr_2_LC_16_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31583),
            .lcout(\PWMInstance3.PWMPulseWidthCountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38636),
            .ce(N__29308),
            .sr(N__35784));
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_16_13_4 .C_ON=1'b0;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_16_13_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_16_13_4 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \PWMInstance3.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_16_13_4  (
            .in0(N__29133),
            .in1(N__29127),
            .in2(N__29175),
            .in3(N__29152),
            .lcout(\PWMInstance3.un1_PWMPulseWidthCount_0_I_21_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance3.PWMPulseWidthCount_esr_14_LC_16_13_5 .C_ON=1'b0;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_14_LC_16_13_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_14_LC_16_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance3.PWMPulseWidthCount_esr_14_LC_16_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34401),
            .lcout(\PWMInstance3.PWMPulseWidthCountZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38636),
            .ce(N__29308),
            .sr(N__35784));
    defparam \PWMInstance3.PWMPulseWidthCount_esr_15_LC_16_13_6 .C_ON=1'b0;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_15_LC_16_13_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_15_LC_16_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance3.PWMPulseWidthCount_esr_15_LC_16_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31903),
            .lcout(\PWMInstance3.PWMPulseWidthCountZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38636),
            .ce(N__29308),
            .sr(N__35784));
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_16_13_7 .C_ON=1'b0;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_16_13_7 .SEQ_MODE=4'b0000;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_16_13_7 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance3.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_16_13_7  (
            .in0(N__29121),
            .in1(N__29115),
            .in2(N__29088),
            .in3(N__29107),
            .lcout(\PWMInstance3.un1_PWMPulseWidthCount_0_I_39_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance3.periodCounter_RNIMJ9L_0_LC_16_14_0 .C_ON=1'b0;
    defparam \PWMInstance3.periodCounter_RNIMJ9L_0_LC_16_14_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance3.periodCounter_RNIMJ9L_0_LC_16_14_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \PWMInstance3.periodCounter_RNIMJ9L_0_LC_16_14_0  (
            .in0(N__29054),
            .in1(N__29083),
            .in2(N__29262),
            .in3(N__29479),
            .lcout(\PWMInstance3.un1_periodCounter12_1_0_a2_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_16_14_1 .C_ON=1'b0;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_16_14_1 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance3.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_16_14_1  (
            .in0(N__29013),
            .in1(N__29053),
            .in2(N__29040),
            .in3(N__29019),
            .lcout(\PWMInstance3.un1_PWMPulseWidthCount_0_I_1_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance3.PWMPulseWidthCount_esr_0_LC_16_14_2 .C_ON=1'b0;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_0_LC_16_14_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_0_LC_16_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance3.PWMPulseWidthCount_esr_0_LC_16_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31412),
            .lcout(\PWMInstance3.PWMPulseWidthCountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38623),
            .ce(N__29318),
            .sr(N__35787));
    defparam \PWMInstance3.PWMPulseWidthCount_esr_1_LC_16_14_3 .C_ON=1'b0;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_1_LC_16_14_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_1_LC_16_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance3.PWMPulseWidthCount_esr_1_LC_16_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31280),
            .lcout(\PWMInstance3.PWMPulseWidthCountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38623),
            .ce(N__29318),
            .sr(N__35787));
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_16_14_4 .C_ON=1'b0;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_16_14_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_16_14_4 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance3.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_16_14_4  (
            .in0(N__29325),
            .in1(N__29466),
            .in2(N__29502),
            .in3(N__29480),
            .lcout(\PWMInstance3.un1_PWMPulseWidthCount_0_I_27_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance3.PWMPulseWidthCount_esr_6_LC_16_14_5 .C_ON=1'b0;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_6_LC_16_14_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_6_LC_16_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance3.PWMPulseWidthCount_esr_6_LC_16_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31094),
            .lcout(\PWMInstance3.PWMPulseWidthCountZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38623),
            .ce(N__29318),
            .sr(N__35787));
    defparam \PWMInstance3.PWMPulseWidthCount_esr_7_LC_16_14_6 .C_ON=1'b0;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_7_LC_16_14_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.PWMPulseWidthCount_esr_7_LC_16_14_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \PWMInstance3.PWMPulseWidthCount_esr_7_LC_16_14_6  (
            .in0(N__29413),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PWMInstance3.PWMPulseWidthCountZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38623),
            .ce(N__29318),
            .sr(N__35787));
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_16_14_7 .C_ON=1'b0;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_16_14_7 .SEQ_MODE=4'b0000;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_16_14_7 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \PWMInstance3.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_16_14_7  (
            .in0(N__29274),
            .in1(N__29257),
            .in2(N__29244),
            .in3(N__29223),
            .lcout(\PWMInstance3.un1_PWMPulseWidthCount_0_I_45_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_1_c_LC_16_15_0 .C_ON=1'b1;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_1_c_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_1_c_LC_16_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance3.un1_PWMPulseWidthCount_0_I_1_c_LC_16_15_0  (
            .in0(_gnd_net_),
            .in1(N__29214),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_15_0_),
            .carryout(\PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_9_c_LC_16_15_1 .C_ON=1'b1;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_9_c_LC_16_15_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_9_c_LC_16_15_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance3.un1_PWMPulseWidthCount_0_I_9_c_LC_16_15_1  (
            .in0(_gnd_net_),
            .in1(N__29208),
            .in2(N__32579),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_0 ),
            .carryout(\PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_15_c_LC_16_15_2 .C_ON=1'b1;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_15_c_LC_16_15_2 .SEQ_MODE=4'b0000;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_15_c_LC_16_15_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance3.un1_PWMPulseWidthCount_0_I_15_c_LC_16_15_2  (
            .in0(_gnd_net_),
            .in1(N__29199),
            .in2(N__32573),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_1 ),
            .carryout(\PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_27_c_LC_16_15_3 .C_ON=1'b1;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_27_c_LC_16_15_3 .SEQ_MODE=4'b0000;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_27_c_LC_16_15_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance3.un1_PWMPulseWidthCount_0_I_27_c_LC_16_15_3  (
            .in0(_gnd_net_),
            .in1(N__29187),
            .in2(N__32577),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_2 ),
            .carryout(\PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_45_c_LC_16_15_4 .C_ON=1'b1;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_45_c_LC_16_15_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_45_c_LC_16_15_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance3.un1_PWMPulseWidthCount_0_I_45_c_LC_16_15_4  (
            .in0(_gnd_net_),
            .in1(N__29820),
            .in2(N__32575),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_3 ),
            .carryout(\PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_33_c_LC_16_15_5 .C_ON=1'b1;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_33_c_LC_16_15_5 .SEQ_MODE=4'b0000;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_33_c_LC_16_15_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance3.un1_PWMPulseWidthCount_0_I_33_c_LC_16_15_5  (
            .in0(_gnd_net_),
            .in1(N__29814),
            .in2(N__32578),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_4 ),
            .carryout(\PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_39_c_LC_16_15_6 .C_ON=1'b1;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_39_c_LC_16_15_6 .SEQ_MODE=4'b0000;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_39_c_LC_16_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance3.un1_PWMPulseWidthCount_0_I_39_c_LC_16_15_6  (
            .in0(_gnd_net_),
            .in1(N__29805),
            .in2(N__32574),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_5 ),
            .carryout(\PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_21_c_LC_16_15_7 .C_ON=1'b1;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_21_c_LC_16_15_7 .SEQ_MODE=4'b0000;
    defparam \PWMInstance3.un1_PWMPulseWidthCount_0_I_21_c_LC_16_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance3.un1_PWMPulseWidthCount_0_I_21_c_LC_16_15_7  (
            .in0(_gnd_net_),
            .in1(N__29796),
            .in2(N__32576),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_6 ),
            .carryout(\PWMInstance3.un1_PWMPulseWidthCount_0_data_tmp_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance3.out_LC_16_16_0 .C_ON=1'b0;
    defparam \PWMInstance3.out_LC_16_16_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance3.out_LC_16_16_0 .LUT_INIT=16'b1111101011110010;
    LogicCell40 \PWMInstance3.out_LC_16_16_0  (
            .in0(N__29717),
            .in1(N__29787),
            .in2(N__29775),
            .in3(N__29730),
            .lcout(PWM3_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38602),
            .ce(),
            .sr(N__35794));
    defparam \QuadInstance7.delayedCh_A_0_LC_16_18_2 .C_ON=1'b0;
    defparam \QuadInstance7.delayedCh_A_0_LC_16_18_2 .SEQ_MODE=4'b1000;
    defparam \QuadInstance7.delayedCh_A_0_LC_16_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance7.delayedCh_A_0_LC_16_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29706),
            .lcout(\QuadInstance7.delayedCh_AZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38584),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_5_LC_17_3_6 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_5_LC_17_3_6 .SEQ_MODE=4'b1000;
    defparam \QuadInstance0.Quad_5_LC_17_3_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance0.Quad_5_LC_17_3_6  (
            .in0(N__36346),
            .in1(N__33109),
            .in2(_gnd_net_),
            .in3(N__29832),
            .lcout(dataRead0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38722),
            .ce(),
            .sr(N__35725));
    defparam \QuadInstance4.Quad_10_LC_17_4_0 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_10_LC_17_4_0 .SEQ_MODE=4'b1000;
    defparam \QuadInstance4.Quad_10_LC_17_4_0 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \QuadInstance4.Quad_10_LC_17_4_0  (
            .in0(N__36165),
            .in1(_gnd_net_),
            .in2(N__29676),
            .in3(N__29661),
            .lcout(dataRead4_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38719),
            .ce(),
            .sr(N__35735));
    defparam \QuadInstance4.Quad_14_LC_17_4_2 .C_ON=1'b0;
    defparam \QuadInstance4.Quad_14_LC_17_4_2 .SEQ_MODE=4'b1000;
    defparam \QuadInstance4.Quad_14_LC_17_4_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \QuadInstance4.Quad_14_LC_17_4_2  (
            .in0(N__34416),
            .in1(N__29660),
            .in2(_gnd_net_),
            .in3(N__29979),
            .lcout(dataRead4_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38719),
            .ce(),
            .sr(N__35735));
    defparam \QuadInstance0.delayedCh_B_1_LC_17_5_1 .C_ON=1'b0;
    defparam \QuadInstance0.delayedCh_B_1_LC_17_5_1 .SEQ_MODE=4'b1000;
    defparam \QuadInstance0.delayedCh_B_1_LC_17_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance0.delayedCh_B_1_LC_17_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29934),
            .lcout(\QuadInstance0.delayedCh_BZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38712),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance4.delayedCh_B_1_LC_17_5_7 .C_ON=1'b0;
    defparam \QuadInstance4.delayedCh_B_1_LC_17_5_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance4.delayedCh_B_1_LC_17_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance4.delayedCh_B_1_LC_17_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29919),
            .lcout(\QuadInstance4.delayedCh_BZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38712),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.un1_Quad_cry_0_c_LC_17_6_0 .C_ON=1'b1;
    defparam \QuadInstance0.un1_Quad_cry_0_c_LC_17_6_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.un1_Quad_cry_0_c_LC_17_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \QuadInstance0.un1_Quad_cry_0_c_LC_17_6_0  (
            .in0(_gnd_net_),
            .in1(N__34046),
            .in2(N__30317),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_6_0_),
            .carryout(\QuadInstance0.un1_Quad_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_RNO_0_1_LC_17_6_1 .C_ON=1'b1;
    defparam \QuadInstance0.Quad_RNO_0_1_LC_17_6_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNO_0_1_LC_17_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance0.Quad_RNO_0_1_LC_17_6_1  (
            .in0(_gnd_net_),
            .in1(N__32729),
            .in2(N__32697),
            .in3(N__29880),
            .lcout(\QuadInstance0.Quad_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\QuadInstance0.un1_Quad_cry_0 ),
            .carryout(\QuadInstance0.un1_Quad_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_RNO_0_2_LC_17_6_2 .C_ON=1'b1;
    defparam \QuadInstance0.Quad_RNO_0_2_LC_17_6_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNO_0_2_LC_17_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance0.Quad_RNO_0_2_LC_17_6_2  (
            .in0(_gnd_net_),
            .in1(N__32657),
            .in2(N__32637),
            .in3(N__29868),
            .lcout(\QuadInstance0.Quad_RNO_0_0_2 ),
            .ltout(),
            .carryin(\QuadInstance0.un1_Quad_cry_1 ),
            .carryout(\QuadInstance0.un1_Quad_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_RNO_0_3_LC_17_6_3 .C_ON=1'b1;
    defparam \QuadInstance0.Quad_RNO_0_3_LC_17_6_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNO_0_3_LC_17_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance0.Quad_RNO_0_3_LC_17_6_3  (
            .in0(_gnd_net_),
            .in1(N__34176),
            .in2(N__34218),
            .in3(N__29850),
            .lcout(\QuadInstance0.Quad_RNO_0_0_3 ),
            .ltout(),
            .carryin(\QuadInstance0.un1_Quad_cry_2 ),
            .carryout(\QuadInstance0.un1_Quad_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_RNO_0_4_LC_17_6_4 .C_ON=1'b1;
    defparam \QuadInstance0.Quad_RNO_0_4_LC_17_6_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNO_0_4_LC_17_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance0.Quad_RNO_0_4_LC_17_6_4  (
            .in0(_gnd_net_),
            .in1(N__34163),
            .in2(N__34134),
            .in3(N__29835),
            .lcout(\QuadInstance0.Quad_RNO_0_0_4 ),
            .ltout(),
            .carryin(\QuadInstance0.un1_Quad_cry_3 ),
            .carryout(\QuadInstance0.un1_Quad_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_RNO_0_5_LC_17_6_5 .C_ON=1'b1;
    defparam \QuadInstance0.Quad_RNO_0_5_LC_17_6_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNO_0_5_LC_17_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance0.Quad_RNO_0_5_LC_17_6_5  (
            .in0(_gnd_net_),
            .in1(N__34121),
            .in2(N__34098),
            .in3(N__29823),
            .lcout(\QuadInstance0.Quad_RNO_0_0_5 ),
            .ltout(),
            .carryin(\QuadInstance0.un1_Quad_cry_4 ),
            .carryout(\QuadInstance0.un1_Quad_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_RNO_0_6_LC_17_6_6 .C_ON=1'b1;
    defparam \QuadInstance0.Quad_RNO_0_6_LC_17_6_6 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNO_0_6_LC_17_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance0.Quad_RNO_0_6_LC_17_6_6  (
            .in0(_gnd_net_),
            .in1(N__33980),
            .in2(N__33867),
            .in3(N__30231),
            .lcout(\QuadInstance0.Quad_RNO_0_0_6 ),
            .ltout(),
            .carryin(\QuadInstance0.un1_Quad_cry_5 ),
            .carryout(\QuadInstance0.un1_Quad_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_RNO_0_7_LC_17_6_7 .C_ON=1'b1;
    defparam \QuadInstance0.Quad_RNO_0_7_LC_17_6_7 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNO_0_7_LC_17_6_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance0.Quad_RNO_0_7_LC_17_6_7  (
            .in0(_gnd_net_),
            .in1(N__30228),
            .in2(N__30213),
            .in3(N__30198),
            .lcout(\QuadInstance0.Quad_RNO_0_0_7 ),
            .ltout(),
            .carryin(\QuadInstance0.un1_Quad_cry_6 ),
            .carryout(\QuadInstance0.un1_Quad_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_RNO_0_8_LC_17_7_0 .C_ON=1'b1;
    defparam \QuadInstance0.Quad_RNO_0_8_LC_17_7_0 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNO_0_8_LC_17_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance0.Quad_RNO_0_8_LC_17_7_0  (
            .in0(_gnd_net_),
            .in1(N__30195),
            .in2(N__30180),
            .in3(N__30165),
            .lcout(\QuadInstance0.Quad_RNO_0_0_8 ),
            .ltout(),
            .carryin(bfn_17_7_0_),
            .carryout(\QuadInstance0.un1_Quad_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_RNO_0_9_LC_17_7_1 .C_ON=1'b1;
    defparam \QuadInstance0.Quad_RNO_0_9_LC_17_7_1 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNO_0_9_LC_17_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance0.Quad_RNO_0_9_LC_17_7_1  (
            .in0(_gnd_net_),
            .in1(N__30162),
            .in2(N__30129),
            .in3(N__30105),
            .lcout(\QuadInstance0.Quad_RNO_0_0_9 ),
            .ltout(),
            .carryin(\QuadInstance0.un1_Quad_cry_8 ),
            .carryout(\QuadInstance0.un1_Quad_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_RNO_0_10_LC_17_7_2 .C_ON=1'b1;
    defparam \QuadInstance0.Quad_RNO_0_10_LC_17_7_2 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNO_0_10_LC_17_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance0.Quad_RNO_0_10_LC_17_7_2  (
            .in0(_gnd_net_),
            .in1(N__32687),
            .in2(N__32670),
            .in3(N__30102),
            .lcout(\QuadInstance0.Quad_RNO_0_0_10 ),
            .ltout(),
            .carryin(\QuadInstance0.un1_Quad_cry_9 ),
            .carryout(\QuadInstance0.un1_Quad_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_RNO_0_11_LC_17_7_3 .C_ON=1'b1;
    defparam \QuadInstance0.Quad_RNO_0_11_LC_17_7_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNO_0_11_LC_17_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance0.Quad_RNO_0_11_LC_17_7_3  (
            .in0(_gnd_net_),
            .in1(N__30098),
            .in2(N__30075),
            .in3(N__30057),
            .lcout(\QuadInstance0.Quad_RNO_0_0_11 ),
            .ltout(),
            .carryin(\QuadInstance0.un1_Quad_cry_10 ),
            .carryout(\QuadInstance0.un1_Quad_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_RNO_0_12_LC_17_7_4 .C_ON=1'b1;
    defparam \QuadInstance0.Quad_RNO_0_12_LC_17_7_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNO_0_12_LC_17_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance0.Quad_RNO_0_12_LC_17_7_4  (
            .in0(_gnd_net_),
            .in1(N__30054),
            .in2(N__30033),
            .in3(N__30018),
            .lcout(\QuadInstance0.Quad_RNO_0_0_12 ),
            .ltout(),
            .carryin(\QuadInstance0.un1_Quad_cry_11 ),
            .carryout(\QuadInstance0.un1_Quad_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_RNO_0_13_LC_17_7_5 .C_ON=1'b1;
    defparam \QuadInstance0.Quad_RNO_0_13_LC_17_7_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNO_0_13_LC_17_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance0.Quad_RNO_0_13_LC_17_7_5  (
            .in0(_gnd_net_),
            .in1(N__30014),
            .in2(N__29997),
            .in3(N__29982),
            .lcout(\QuadInstance0.Quad_RNO_0_0_13 ),
            .ltout(),
            .carryin(\QuadInstance0.un1_Quad_cry_12 ),
            .carryout(\QuadInstance0.un1_Quad_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_RNO_0_14_LC_17_7_6 .C_ON=1'b1;
    defparam \QuadInstance0.Quad_RNO_0_14_LC_17_7_6 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNO_0_14_LC_17_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \QuadInstance0.Quad_RNO_0_14_LC_17_7_6  (
            .in0(_gnd_net_),
            .in1(N__34224),
            .in2(N__34250),
            .in3(N__30597),
            .lcout(\QuadInstance0.Quad_RNO_0_0_14 ),
            .ltout(),
            .carryin(\QuadInstance0.un1_Quad_cry_13 ),
            .carryout(\QuadInstance0.un1_Quad_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_15_LC_17_7_7 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_15_LC_17_7_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance0.Quad_15_LC_17_7_7 .LUT_INIT=16'b1101000111100010;
    LogicCell40 \QuadInstance0.Quad_15_LC_17_7_7  (
            .in0(N__30594),
            .in1(N__33044),
            .in2(N__31917),
            .in3(N__30585),
            .lcout(dataRead0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38699),
            .ce(),
            .sr(N__35753));
    defparam OutReg_esr_RNO_2_2_LC_17_8_0.C_ON=1'b0;
    defparam OutReg_esr_RNO_2_2_LC_17_8_0.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_2_2_LC_17_8_0.LUT_INIT=16'b1000100011110011;
    LogicCell40 OutReg_esr_RNO_2_2_LC_17_8_0 (
            .in0(N__30570),
            .in1(N__38154),
            .in2(N__30534),
            .in3(N__30492),
            .lcout(),
            .ltout(OutReg_esr_RNO_2Z0Z_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_esr_RNO_0_2_LC_17_8_1.C_ON=1'b0;
    defparam OutReg_esr_RNO_0_2_LC_17_8_1.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_0_2_LC_17_8_1.LUT_INIT=16'b1111110000110000;
    LogicCell40 OutReg_esr_RNO_0_2_LC_17_8_1 (
            .in0(_gnd_net_),
            .in1(N__37557),
            .in2(N__30480),
            .in3(N__30324),
            .lcout(),
            .ltout(OutReg_esr_RNO_0Z0Z_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_esr_2_LC_17_8_2.C_ON=1'b0;
    defparam OutReg_esr_2_LC_17_8_2.SEQ_MODE=4'b1000;
    defparam OutReg_esr_2_LC_17_8_2.LUT_INIT=16'b1100110011011000;
    LogicCell40 OutReg_esr_2_LC_17_8_2 (
            .in0(N__37332),
            .in1(N__30717),
            .in2(N__30477),
            .in3(N__38932),
            .lcout(OutRegZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38693),
            .ce(N__37224),
            .sr(N__37115));
    defparam OutReg_esr_RNO_3_2_LC_17_8_3.C_ON=1'b0;
    defparam OutReg_esr_RNO_3_2_LC_17_8_3.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_3_2_LC_17_8_3.LUT_INIT=16'b0000001111011101;
    LogicCell40 OutReg_esr_RNO_3_2_LC_17_8_3 (
            .in0(N__30460),
            .in1(N__34885),
            .in2(N__30426),
            .in3(N__34764),
            .lcout(),
            .ltout(OutReg_0_4_i_m3_ns_1_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_esr_RNO_1_2_LC_17_8_4.C_ON=1'b0;
    defparam OutReg_esr_RNO_1_2_LC_17_8_4.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_1_2_LC_17_8_4.LUT_INIT=16'b1100101000001111;
    LogicCell40 OutReg_esr_RNO_1_2_LC_17_8_4 (
            .in0(N__30387),
            .in1(N__30353),
            .in2(N__30327),
            .in3(N__32831),
            .lcout(OutReg_esr_RNO_1Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_4_0_LC_17_9_0.C_ON=1'b0;
    defparam OutReg_ess_RNO_4_0_LC_17_9_0.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_4_0_LC_17_9_0.LUT_INIT=16'b0101010100011011;
    LogicCell40 OutReg_ess_RNO_4_0_LC_17_9_0 (
            .in0(N__37763),
            .in1(N__30318),
            .in2(N__30285),
            .in3(N__38155),
            .lcout(),
            .ltout(OutReg_0_5_i_m3_ns_1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_1_0_LC_17_9_1.C_ON=1'b0;
    defparam OutReg_ess_RNO_1_0_LC_17_9_1.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_1_0_LC_17_9_1.LUT_INIT=16'b1000111110000101;
    LogicCell40 OutReg_ess_RNO_1_0_LC_17_9_1 (
            .in0(N__38156),
            .in1(N__30951),
            .in2(N__30918),
            .in3(N__30915),
            .lcout(),
            .ltout(OutReg_ess_RNO_1Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_0_LC_17_9_2.C_ON=1'b0;
    defparam OutReg_ess_0_LC_17_9_2.SEQ_MODE=4'b1001;
    defparam OutReg_ess_0_LC_17_9_2.LUT_INIT=16'b1000100011000000;
    LogicCell40 OutReg_ess_0_LC_17_9_2 (
            .in0(N__30747),
            .in1(N__34944),
            .in2(N__30885),
            .in3(N__37562),
            .lcout(OutRegZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38685),
            .ce(N__37210),
            .sr(N__37128));
    defparam OutReg_ess_RNO_3_0_LC_17_9_3.C_ON=1'b0;
    defparam OutReg_ess_RNO_3_0_LC_17_9_3.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_3_0_LC_17_9_3.LUT_INIT=16'b0001000111001111;
    LogicCell40 OutReg_ess_RNO_3_0_LC_17_9_3 (
            .in0(N__30882),
            .in1(N__37761),
            .in2(N__30849),
            .in3(N__32949),
            .lcout(),
            .ltout(OutReg_0_4_i_m3_ns_1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_0_0_LC_17_9_4.C_ON=1'b0;
    defparam OutReg_ess_RNO_0_0_LC_17_9_4.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_0_0_LC_17_9_4.LUT_INIT=16'b1000111110000101;
    LogicCell40 OutReg_ess_RNO_0_0_LC_17_9_4 (
            .in0(N__37762),
            .in1(N__30809),
            .in2(N__30780),
            .in3(N__30777),
            .lcout(OutReg_ess_RNO_0Z0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_1_LC_17_9_6.C_ON=1'b0;
    defparam OutReg_ess_1_LC_17_9_6.SEQ_MODE=4'b1001;
    defparam OutReg_ess_1_LC_17_9_6.LUT_INIT=16'b1111000111100000;
    LogicCell40 OutReg_ess_1_LC_17_9_6 (
            .in0(N__37323),
            .in1(N__38913),
            .in2(N__30741),
            .in3(N__30729),
            .lcout(OutRegZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38685),
            .ce(N__37210),
            .sr(N__37128));
    defparam OutReg_esr_RNO_3_8_LC_17_10_1.C_ON=1'b0;
    defparam OutReg_esr_RNO_3_8_LC_17_10_1.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_3_8_LC_17_10_1.LUT_INIT=16'b0000001111011101;
    LogicCell40 OutReg_esr_RNO_3_8_LC_17_10_1 (
            .in0(N__30710),
            .in1(N__34894),
            .in2(N__30675),
            .in3(N__34771),
            .lcout(OutReg_0_4_i_m3_ns_1_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_received_esr_RNI7L871_3_LC_17_10_3.C_ON=1'b0;
    defparam data_received_esr_RNI7L871_3_LC_17_10_3.SEQ_MODE=4'b0000;
    defparam data_received_esr_RNI7L871_3_LC_17_10_3.LUT_INIT=16'b1111111100000001;
    LogicCell40 data_received_esr_RNI7L871_3_LC_17_10_3 (
            .in0(N__37313),
            .in1(N__38878),
            .in2(N__30642),
            .in3(N__39078),
            .lcout(),
            .ltout(data_received_esr_RNI7L871Z0Z_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_received_esr_RNIKE1M2_3_LC_17_10_4.C_ON=1'b0;
    defparam data_received_esr_RNIKE1M2_3_LC_17_10_4.SEQ_MODE=4'b0000;
    defparam data_received_esr_RNIKE1M2_3_LC_17_10_4.LUT_INIT=16'b1111111111110000;
    LogicCell40 data_received_esr_RNIKE1M2_3_LC_17_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30600),
            .in3(N__37060),
            .lcout(N_863_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_received_esr_RNIDPOE1_3_LC_17_10_6.C_ON=1'b0;
    defparam data_received_esr_RNIDPOE1_3_LC_17_10_6.SEQ_MODE=4'b0000;
    defparam data_received_esr_RNIDPOE1_3_LC_17_10_6.LUT_INIT=16'b0001000100000000;
    LogicCell40 data_received_esr_RNIDPOE1_3_LC_17_10_6 (
            .in0(N__38877),
            .in1(N__37312),
            .in2(_gnd_net_),
            .in3(N__31446),
            .lcout(OutReg_0_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.periodCounter_RNIIEMR_13_LC_17_11_0 .C_ON=1'b0;
    defparam \PWMInstance2.periodCounter_RNIIEMR_13_LC_17_11_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance2.periodCounter_RNIIEMR_13_LC_17_11_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \PWMInstance2.periodCounter_RNIIEMR_13_LC_17_11_0  (
            .in0(N__34550),
            .in1(N__35422),
            .in2(N__35154),
            .in3(N__35107),
            .lcout(\PWMInstance2.un1_periodCounter12_1_0_a2_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_17_11_1 .C_ON=1'b0;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_17_11_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_17_11_1 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance2.un1_PWMPulseWidthCount_0_I_1_c_RNO_LC_17_11_1  (
            .in0(N__31137),
            .in1(N__34549),
            .in2(N__35208),
            .in3(N__31287),
            .lcout(\PWMInstance2.un1_PWMPulseWidthCount_0_I_1_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.PWMPulseWidthCount_esr_0_LC_17_11_2 .C_ON=1'b0;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_0_LC_17_11_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_0_LC_17_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance2.PWMPulseWidthCount_esr_0_LC_17_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31437),
            .lcout(\PWMInstance2.PWMPulseWidthCountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38668),
            .ce(N__35861),
            .sr(N__35777));
    defparam \PWMInstance2.PWMPulseWidthCount_esr_1_LC_17_11_3 .C_ON=1'b0;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_1_LC_17_11_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_1_LC_17_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance2.PWMPulseWidthCount_esr_1_LC_17_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31240),
            .lcout(\PWMInstance2.PWMPulseWidthCountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38668),
            .ce(N__35861),
            .sr(N__35777));
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_17_11_4 .C_ON=1'b0;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_17_11_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_17_11_4 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \PWMInstance2.un1_PWMPulseWidthCount_0_I_27_c_RNO_LC_17_11_4  (
            .in0(N__31131),
            .in1(N__30969),
            .in2(N__35153),
            .in3(N__35129),
            .lcout(\PWMInstance2.un1_PWMPulseWidthCount_0_I_27_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.PWMPulseWidthCount_esr_6_LC_17_11_5 .C_ON=1'b0;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_6_LC_17_11_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_6_LC_17_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance2.PWMPulseWidthCount_esr_6_LC_17_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31063),
            .lcout(\PWMInstance2.PWMPulseWidthCountZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38668),
            .ce(N__35861),
            .sr(N__35777));
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_17_11_7 .C_ON=1'b0;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_17_11_7 .SEQ_MODE=4'b0000;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_17_11_7 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance2.un1_PWMPulseWidthCount_0_I_45_c_RNO_LC_17_11_7  (
            .in0(N__30963),
            .in1(N__35455),
            .in2(N__35109),
            .in3(N__30957),
            .lcout(\PWMInstance2.un1_PWMPulseWidthCount_0_I_45_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.out_RNO_0_LC_17_12_0 .C_ON=1'b0;
    defparam \PWMInstance2.out_RNO_0_LC_17_12_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance2.out_RNO_0_LC_17_12_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \PWMInstance2.out_RNO_0_LC_17_12_0  (
            .in0(N__31677),
            .in1(N__31657),
            .in2(N__35334),
            .in3(N__31642),
            .lcout(\PWMInstance2.un1_periodCounter12_1_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.clkCount_0_LC_17_12_1 .C_ON=1'b0;
    defparam \PWMInstance2.clkCount_0_LC_17_12_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.clkCount_0_LC_17_12_1 .LUT_INIT=16'b1010101000000101;
    LogicCell40 \PWMInstance2.clkCount_0_LC_17_12_1  (
            .in0(N__31643),
            .in1(_gnd_net_),
            .in2(N__31664),
            .in3(N__31691),
            .lcout(\PWMInstance2.clkCountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38656),
            .ce(),
            .sr(N__35785));
    defparam \PWMInstance2.PWMPulseWidthCount_esr_ctle_15_LC_17_12_2 .C_ON=1'b0;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_ctle_15_LC_17_12_2 .SEQ_MODE=4'b0000;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_ctle_15_LC_17_12_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \PWMInstance2.PWMPulseWidthCount_esr_ctle_15_LC_17_12_2  (
            .in0(N__31690),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35831),
            .lcout(\PWMInstance2.pwmWrite_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.clkCount_1_LC_17_12_3 .C_ON=1'b0;
    defparam \PWMInstance2.clkCount_1_LC_17_12_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.clkCount_1_LC_17_12_3 .LUT_INIT=16'b1111000000001010;
    LogicCell40 \PWMInstance2.clkCount_1_LC_17_12_3  (
            .in0(N__31644),
            .in1(_gnd_net_),
            .in2(N__31665),
            .in3(N__31692),
            .lcout(\PWMInstance2.clkCountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38656),
            .ce(),
            .sr(N__35785));
    defparam \PWMInstance2.clkCount_RNIV7AK_0_LC_17_12_4 .C_ON=1'b0;
    defparam \PWMInstance2.clkCount_RNIV7AK_0_LC_17_12_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance2.clkCount_RNIV7AK_0_LC_17_12_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \PWMInstance2.clkCount_RNIV7AK_0_LC_17_12_4  (
            .in0(N__31676),
            .in1(N__31656),
            .in2(_gnd_net_),
            .in3(N__31641),
            .lcout(\PWMInstance2.periodCounter12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.periodCounter_RNI6H1B_16_LC_17_12_5 .C_ON=1'b0;
    defparam \PWMInstance2.periodCounter_RNI6H1B_16_LC_17_12_5 .SEQ_MODE=4'b0000;
    defparam \PWMInstance2.periodCounter_RNI6H1B_16_LC_17_12_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \PWMInstance2.periodCounter_RNI6H1B_16_LC_17_12_5  (
            .in0(_gnd_net_),
            .in1(N__35329),
            .in2(_gnd_net_),
            .in3(N__35128),
            .lcout(),
            .ltout(\PWMInstance2.un1_periodCounter12_1_0_a2_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.periodCounter_RNI43DA1_15_LC_17_12_6 .C_ON=1'b0;
    defparam \PWMInstance2.periodCounter_RNI43DA1_15_LC_17_12_6 .SEQ_MODE=4'b0000;
    defparam \PWMInstance2.periodCounter_RNI43DA1_15_LC_17_12_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \PWMInstance2.periodCounter_RNI43DA1_15_LC_17_12_6  (
            .in0(N__35395),
            .in1(N__35206),
            .in2(N__31629),
            .in3(N__34567),
            .lcout(),
            .ltout(\PWMInstance2.un1_periodCounter12_1_0_a2_0_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.periodCounter_RNICCJQ3_10_LC_17_12_7 .C_ON=1'b0;
    defparam \PWMInstance2.periodCounter_RNICCJQ3_10_LC_17_12_7 .SEQ_MODE=4'b0000;
    defparam \PWMInstance2.periodCounter_RNICCJQ3_10_LC_17_12_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \PWMInstance2.periodCounter_RNICCJQ3_10_LC_17_12_7  (
            .in0(N__36534),
            .in1(N__31626),
            .in2(N__31620),
            .in3(N__31617),
            .lcout(\PWMInstance2.out_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.periodCounter_RNIJFMR_11_LC_17_13_0 .C_ON=1'b0;
    defparam \PWMInstance2.periodCounter_RNIJFMR_11_LC_17_13_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance2.periodCounter_RNIJFMR_11_LC_17_13_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \PWMInstance2.periodCounter_RNIJFMR_11_LC_17_13_0  (
            .in0(N__35180),
            .in1(N__35456),
            .in2(N__36200),
            .in3(N__35237),
            .lcout(\PWMInstance2.un1_periodCounter12_1_0_a2_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_17_13_1 .C_ON=1'b0;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_17_13_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_17_13_1 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \PWMInstance2.un1_PWMPulseWidthCount_0_I_9_c_RNO_LC_17_13_1  (
            .in0(N__31935),
            .in1(N__35181),
            .in2(N__31455),
            .in3(N__36597),
            .lcout(\PWMInstance2.un1_PWMPulseWidthCount_0_I_9_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.PWMPulseWidthCount_esr_2_LC_17_13_2 .C_ON=1'b0;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_2_LC_17_13_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_2_LC_17_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance2.PWMPulseWidthCount_esr_2_LC_17_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31584),
            .lcout(\PWMInstance2.PWMPulseWidthCountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38646),
            .ce(N__35853),
            .sr(N__35788));
    defparam \PWMInstance2.PWMPulseWidthCount_esr_3_LC_17_13_3 .C_ON=1'b0;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_3_LC_17_13_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_3_LC_17_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance2.PWMPulseWidthCount_esr_3_LC_17_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32033),
            .lcout(\PWMInstance2.PWMPulseWidthCountZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38646),
            .ce(N__35853),
            .sr(N__35788));
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_17_13_4 .C_ON=1'b0;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_17_13_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_17_13_4 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance2.un1_PWMPulseWidthCount_0_I_21_c_RNO_LC_17_13_4  (
            .in0(N__31737),
            .in1(N__31929),
            .in2(N__35400),
            .in3(N__36616),
            .lcout(\PWMInstance2.un1_PWMPulseWidthCount_0_I_21_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.PWMPulseWidthCount_esr_14_LC_17_13_5 .C_ON=1'b0;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_14_LC_17_13_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_14_LC_17_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance2.PWMPulseWidthCount_esr_14_LC_17_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34400),
            .lcout(\PWMInstance2.PWMPulseWidthCountZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38646),
            .ce(N__35853),
            .sr(N__35788));
    defparam \PWMInstance2.PWMPulseWidthCount_esr_15_LC_17_13_6 .C_ON=1'b0;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_15_LC_17_13_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_15_LC_17_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance2.PWMPulseWidthCount_esr_15_LC_17_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31904),
            .lcout(\PWMInstance2.PWMPulseWidthCountZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38646),
            .ce(N__35853),
            .sr(N__35788));
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_17_13_7 .C_ON=1'b0;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_17_13_7 .SEQ_MODE=4'b0000;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_17_13_7 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \PWMInstance2.un1_PWMPulseWidthCount_0_I_39_c_RNO_LC_17_13_7  (
            .in0(N__31731),
            .in1(N__31719),
            .in2(N__35427),
            .in3(N__36556),
            .lcout(\PWMInstance2.un1_PWMPulseWidthCount_0_I_39_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_1_c_LC_17_14_0 .C_ON=1'b1;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_1_c_LC_17_14_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_1_c_LC_17_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance2.un1_PWMPulseWidthCount_0_I_1_c_LC_17_14_0  (
            .in0(_gnd_net_),
            .in1(N__31710),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_14_0_),
            .carryout(\PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_9_c_LC_17_14_1 .C_ON=1'b1;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_9_c_LC_17_14_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_9_c_LC_17_14_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance2.un1_PWMPulseWidthCount_0_I_9_c_LC_17_14_1  (
            .in0(_gnd_net_),
            .in1(N__32390),
            .in2(N__31701),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_0 ),
            .carryout(\PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_15_c_LC_17_14_2 .C_ON=1'b1;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_15_c_LC_17_14_2 .SEQ_MODE=4'b0000;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_15_c_LC_17_14_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance2.un1_PWMPulseWidthCount_0_I_15_c_LC_17_14_2  (
            .in0(_gnd_net_),
            .in1(N__35214),
            .in2(N__32494),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_1 ),
            .carryout(\PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_27_c_LC_17_14_3 .C_ON=1'b1;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_27_c_LC_17_14_3 .SEQ_MODE=4'b0000;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_27_c_LC_17_14_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance2.un1_PWMPulseWidthCount_0_I_27_c_LC_17_14_3  (
            .in0(_gnd_net_),
            .in1(N__32383),
            .in2(N__32619),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_2 ),
            .carryout(\PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_45_c_LC_17_14_4 .C_ON=1'b1;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_45_c_LC_17_14_4 .SEQ_MODE=4'b0000;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_45_c_LC_17_14_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance2.un1_PWMPulseWidthCount_0_I_45_c_LC_17_14_4  (
            .in0(_gnd_net_),
            .in1(N__32607),
            .in2(N__32496),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_3 ),
            .carryout(\PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_33_c_LC_17_14_5 .C_ON=1'b1;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_33_c_LC_17_14_5 .SEQ_MODE=4'b0000;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_33_c_LC_17_14_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance2.un1_PWMPulseWidthCount_0_I_33_c_LC_17_14_5  (
            .in0(_gnd_net_),
            .in1(N__36174),
            .in2(N__32518),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_4 ),
            .carryout(\PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_39_c_LC_17_14_6 .C_ON=1'b1;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_39_c_LC_17_14_6 .SEQ_MODE=4'b0000;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_39_c_LC_17_14_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance2.un1_PWMPulseWidthCount_0_I_39_c_LC_17_14_6  (
            .in0(_gnd_net_),
            .in1(N__32598),
            .in2(N__32495),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_5 ),
            .carryout(\PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_21_c_LC_17_14_7 .C_ON=1'b1;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_21_c_LC_17_14_7 .SEQ_MODE=4'b0000;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_21_c_LC_17_14_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PWMInstance2.un1_PWMPulseWidthCount_0_I_21_c_LC_17_14_7  (
            .in0(_gnd_net_),
            .in1(N__32382),
            .in2(N__32172),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_6 ),
            .carryout(\PWMInstance2.un1_PWMPulseWidthCount_0_data_tmp_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.out_LC_17_15_0 .C_ON=1'b0;
    defparam \PWMInstance2.out_LC_17_15_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.out_LC_17_15_0 .LUT_INIT=16'b1111101011110010;
    LogicCell40 \PWMInstance2.out_LC_17_15_0  (
            .in0(N__32141),
            .in1(N__32163),
            .in2(N__35376),
            .in3(N__32154),
            .lcout(PWM2_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38624),
            .ce(),
            .sr(N__35795));
    defparam MOSIr_0_LC_18_1_3.C_ON=1'b0;
    defparam MOSIr_0_LC_18_1_3.SEQ_MODE=4'b1000;
    defparam MOSIr_0_LC_18_1_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 MOSIr_0_LC_18_1_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32130),
            .lcout(MOSIrZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38723),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance1.delayedCh_A_0_LC_18_1_7 .C_ON=1'b0;
    defparam \QuadInstance1.delayedCh_A_0_LC_18_1_7 .SEQ_MODE=4'b1000;
    defparam \QuadInstance1.delayedCh_A_0_LC_18_1_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance1.delayedCh_A_0_LC_18_1_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32124),
            .lcout(\QuadInstance1.delayedCh_AZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38723),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.delayedCh_A_1_LC_18_5_0 .C_ON=1'b0;
    defparam \QuadInstance0.delayedCh_A_1_LC_18_5_0 .SEQ_MODE=4'b1000;
    defparam \QuadInstance0.delayedCh_A_1_LC_18_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance0.delayedCh_A_1_LC_18_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32106),
            .lcout(\QuadInstance0.delayedCh_AZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38720),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.delayedCh_A_2_LC_18_5_1 .C_ON=1'b0;
    defparam \QuadInstance0.delayedCh_A_2_LC_18_5_1 .SEQ_MODE=4'b1000;
    defparam \QuadInstance0.delayedCh_A_2_LC_18_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \QuadInstance0.delayedCh_A_2_LC_18_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34534),
            .lcout(\QuadInstance0.delayedCh_AZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38720),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.delayedCh_B_2_LC_18_5_4 .C_ON=1'b0;
    defparam \QuadInstance0.delayedCh_B_2_LC_18_5_4 .SEQ_MODE=4'b1000;
    defparam \QuadInstance0.delayedCh_B_2_LC_18_5_4 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \QuadInstance0.delayedCh_B_2_LC_18_5_4  (
            .in0(_gnd_net_),
            .in1(N__32751),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\QuadInstance0.delayedCh_BZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38720),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_esr_RNO_4_10_LC_18_6_0.C_ON=1'b0;
    defparam OutReg_esr_RNO_4_10_LC_18_6_0.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_4_10_LC_18_6_0.LUT_INIT=16'b0001101000011111;
    LogicCell40 OutReg_esr_RNO_4_10_LC_18_6_0 (
            .in0(N__32944),
            .in1(N__32866),
            .in2(N__32840),
            .in3(N__32683),
            .lcout(OutReg_0_5_i_m3_ns_1_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_10_LC_18_6_1 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_10_LC_18_6_1 .SEQ_MODE=4'b1000;
    defparam \QuadInstance0.Quad_10_LC_18_6_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \QuadInstance0.Quad_10_LC_18_6_1  (
            .in0(N__33048),
            .in1(_gnd_net_),
            .in2(N__36164),
            .in3(N__32757),
            .lcout(dataRead0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38713),
            .ce(),
            .sr(N__35754));
    defparam \QuadInstance0.delayedCh_A_RNICHIP_2_LC_18_6_3 .C_ON=1'b0;
    defparam \QuadInstance0.delayedCh_A_RNICHIP_2_LC_18_6_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.delayedCh_A_RNICHIP_2_LC_18_6_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \QuadInstance0.delayedCh_A_RNICHIP_2_LC_18_6_3  (
            .in0(N__32627),
            .in1(N__32750),
            .in2(N__34536),
            .in3(N__32739),
            .lcout(\QuadInstance0.count_enable ),
            .ltout(\QuadInstance0.count_enable_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_RNIGEBH1_1_LC_18_6_4 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_RNIGEBH1_1_LC_18_6_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNIGEBH1_1_LC_18_6_4 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance0.Quad_RNIGEBH1_1_LC_18_6_4  (
            .in0(N__32733),
            .in1(N__33045),
            .in2(N__32700),
            .in3(N__33903),
            .lcout(\QuadInstance0.Quad_RNIGEBH1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_RNI0L8Q1_10_LC_18_6_5 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_RNI0L8Q1_10_LC_18_6_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNI0L8Q1_10_LC_18_6_5 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \QuadInstance0.Quad_RNI0L8Q1_10_LC_18_6_5  (
            .in0(N__33047),
            .in1(N__33924),
            .in2(N__32688),
            .in3(N__34028),
            .lcout(\QuadInstance0.Quad_RNI0L8Q1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_RNIHFBH1_2_LC_18_6_6 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_RNIHFBH1_2_LC_18_6_6 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNIHFBH1_2_LC_18_6_6 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \QuadInstance0.Quad_RNIHFBH1_2_LC_18_6_6  (
            .in0(N__32661),
            .in1(N__33046),
            .in2(N__34048),
            .in3(N__33904),
            .lcout(\QuadInstance0.Quad_RNIHFBH1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.delayedCh_B_RNIK4UJ_2_LC_18_6_7 .C_ON=1'b0;
    defparam \QuadInstance0.delayedCh_B_RNIK4UJ_2_LC_18_6_7 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.delayedCh_B_RNIK4UJ_2_LC_18_6_7 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \QuadInstance0.delayedCh_B_RNIK4UJ_2_LC_18_6_7  (
            .in0(N__32628),
            .in1(_gnd_net_),
            .in2(N__34535),
            .in3(N__34511),
            .lcout(\QuadInstance0.un1_count_enable_i_a2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_14_LC_18_7_1 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_14_LC_18_7_1 .SEQ_MODE=4'b1000;
    defparam \QuadInstance0.Quad_14_LC_18_7_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \QuadInstance0.Quad_14_LC_18_7_1  (
            .in0(N__34415),
            .in1(_gnd_net_),
            .in2(N__33053),
            .in3(N__34257),
            .lcout(dataRead0_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38707),
            .ce(),
            .sr(N__35758));
    defparam \QuadInstance0.Quad_RNI4P8Q1_14_LC_18_7_3 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_RNI4P8Q1_14_LC_18_7_3 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNI4P8Q1_14_LC_18_7_3 .LUT_INIT=16'b1010001010100010;
    LogicCell40 \QuadInstance0.Quad_RNI4P8Q1_14_LC_18_7_3  (
            .in0(N__34047),
            .in1(N__33913),
            .in2(N__33052),
            .in3(N__34249),
            .lcout(\QuadInstance0.Quad_RNI4P8Q1Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_RNIIGBH1_3_LC_18_7_4 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_RNIIGBH1_3_LC_18_7_4 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNIIGBH1_3_LC_18_7_4 .LUT_INIT=16'b1010101000001010;
    LogicCell40 \QuadInstance0.Quad_RNIIGBH1_3_LC_18_7_4  (
            .in0(N__34030),
            .in1(N__34207),
            .in2(N__33925),
            .in3(N__33012),
            .lcout(\QuadInstance0.Quad_RNIIGBH1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_RNIJHBH1_4_LC_18_7_5 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_RNIJHBH1_4_LC_18_7_5 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNIJHBH1_4_LC_18_7_5 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \QuadInstance0.Quad_RNIJHBH1_4_LC_18_7_5  (
            .in0(N__33014),
            .in1(N__34029),
            .in2(N__34170),
            .in3(N__33905),
            .lcout(\QuadInstance0.Quad_RNIJHBH1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_RNIKIBH1_5_LC_18_7_6 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_RNIKIBH1_5_LC_18_7_6 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNIKIBH1_5_LC_18_7_6 .LUT_INIT=16'b1010101000001010;
    LogicCell40 \QuadInstance0.Quad_RNIKIBH1_5_LC_18_7_6  (
            .in0(N__34032),
            .in1(N__34125),
            .in2(N__33926),
            .in3(N__33013),
            .lcout(\QuadInstance0.Quad_RNIKIBH1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \QuadInstance0.Quad_RNILJBH1_6_LC_18_7_7 .C_ON=1'b0;
    defparam \QuadInstance0.Quad_RNILJBH1_6_LC_18_7_7 .SEQ_MODE=4'b0000;
    defparam \QuadInstance0.Quad_RNILJBH1_6_LC_18_7_7 .LUT_INIT=16'b1000100011001100;
    LogicCell40 \QuadInstance0.Quad_RNILJBH1_6_LC_18_7_7  (
            .in0(N__33015),
            .in1(N__34031),
            .in2(N__33984),
            .in3(N__33909),
            .lcout(\QuadInstance0.Quad_RNILJBH1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam quadWrite_0_LC_18_8_0.C_ON=1'b0;
    defparam quadWrite_0_LC_18_8_0.SEQ_MODE=4'b1000;
    defparam quadWrite_0_LC_18_8_0.LUT_INIT=16'b0001000000000000;
    LogicCell40 quadWrite_0_LC_18_8_0 (
            .in0(N__33851),
            .in1(N__33619),
            .in2(N__33400),
            .in3(N__33232),
            .lcout(quadWriteZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38700),
            .ce(),
            .sr(_gnd_net_));
    defparam MOSIr_1_LC_18_8_1.C_ON=1'b0;
    defparam MOSIr_1_LC_18_8_1.SEQ_MODE=4'b1000;
    defparam MOSIr_1_LC_18_8_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 MOSIr_1_LC_18_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32958),
            .lcout(MOSIrZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38700),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_esr_RNO_2_10_LC_18_8_4.C_ON=1'b0;
    defparam OutReg_esr_RNO_2_10_LC_18_8_4.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_2_10_LC_18_8_4.LUT_INIT=16'b1000100011110011;
    LogicCell40 OutReg_esr_RNO_2_10_LC_18_8_4 (
            .in0(N__35060),
            .in1(N__38159),
            .in2(N__35025),
            .in3(N__34989),
            .lcout(OutReg_esr_RNO_2Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam bit_count_RNI5AMB_0_LC_18_9_2.C_ON=1'b0;
    defparam bit_count_RNI5AMB_0_LC_18_9_2.SEQ_MODE=4'b0000;
    defparam bit_count_RNI5AMB_0_LC_18_9_2.LUT_INIT=16'b1111111111110111;
    LogicCell40 bit_count_RNI5AMB_0_LC_18_9_2 (
            .in0(N__37961),
            .in1(N__37886),
            .in2(N__34980),
            .in3(N__37812),
            .lcout(un1_OutReg51_4_0_i_o3_2),
            .ltout(un1_OutReg51_4_0_i_o3_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_2_0_LC_18_9_3.C_ON=1'b0;
    defparam OutReg_ess_RNO_2_0_LC_18_9_3.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_2_0_LC_18_9_3.LUT_INIT=16'b0000000000001111;
    LogicCell40 OutReg_ess_RNO_2_0_LC_18_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34947),
            .in3(N__38912),
            .lcout(OutReg_21_m_0_a2_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_esr_RNO_0_10_LC_18_9_4.C_ON=1'b0;
    defparam OutReg_esr_RNO_0_10_LC_18_9_4.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_0_10_LC_18_9_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 OutReg_esr_RNO_0_10_LC_18_9_4 (
            .in0(N__37561),
            .in1(N__34578),
            .in2(_gnd_net_),
            .in3(N__34938),
            .lcout(OutReg_esr_RNO_0Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_esr_10_LC_18_10_0.C_ON=1'b0;
    defparam OutReg_esr_10_LC_18_10_0.SEQ_MODE=4'b1000;
    defparam OutReg_esr_10_LC_18_10_0.LUT_INIT=16'b1111000111100000;
    LogicCell40 OutReg_esr_10_LC_18_10_0 (
            .in0(N__38900),
            .in1(N__37322),
            .in2(N__34932),
            .in3(N__34917),
            .lcout(OutRegZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38686),
            .ce(N__37211),
            .sr(N__37099));
    defparam OutReg_esr_RNO_3_10_LC_18_10_1.C_ON=1'b0;
    defparam OutReg_esr_RNO_3_10_LC_18_10_1.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_3_10_LC_18_10_1.LUT_INIT=16'b0001101000011111;
    LogicCell40 OutReg_esr_RNO_3_10_LC_18_10_1 (
            .in0(N__34893),
            .in1(N__34802),
            .in2(N__34773),
            .in3(N__34683),
            .lcout(),
            .ltout(OutReg_0_4_i_m3_ns_1_10_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_esr_RNO_1_10_LC_18_10_2.C_ON=1'b0;
    defparam OutReg_esr_RNO_1_10_LC_18_10_2.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_1_10_LC_18_10_2.LUT_INIT=16'b1100101000001111;
    LogicCell40 OutReg_esr_RNO_1_10_LC_18_10_2 (
            .in0(N__34649),
            .in1(N__34614),
            .in2(N__34581),
            .in3(N__37743),
            .lcout(OutReg_esr_RNO_1Z0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.periodCounter_0_LC_18_11_0 .C_ON=1'b1;
    defparam \PWMInstance2.periodCounter_0_LC_18_11_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.periodCounter_0_LC_18_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance2.periodCounter_0_LC_18_11_0  (
            .in0(_gnd_net_),
            .in1(N__34551),
            .in2(N__34572),
            .in3(N__34571),
            .lcout(\PWMInstance2.periodCounterZ0Z_0 ),
            .ltout(),
            .carryin(bfn_18_11_0_),
            .carryout(\PWMInstance2.un1_periodCounter_2_cry_0 ),
            .clk(N__38677),
            .ce(),
            .sr(N__35310));
    defparam \PWMInstance2.periodCounter_1_LC_18_11_1 .C_ON=1'b1;
    defparam \PWMInstance2.periodCounter_1_LC_18_11_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.periodCounter_1_LC_18_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance2.periodCounter_1_LC_18_11_1  (
            .in0(_gnd_net_),
            .in1(N__35207),
            .in2(_gnd_net_),
            .in3(N__35187),
            .lcout(\PWMInstance2.periodCounterZ0Z_1 ),
            .ltout(),
            .carryin(\PWMInstance2.un1_periodCounter_2_cry_0 ),
            .carryout(\PWMInstance2.un1_periodCounter_2_cry_1 ),
            .clk(N__38677),
            .ce(),
            .sr(N__35310));
    defparam \PWMInstance2.periodCounter_2_LC_18_11_2 .C_ON=1'b1;
    defparam \PWMInstance2.periodCounter_2_LC_18_11_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.periodCounter_2_LC_18_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance2.periodCounter_2_LC_18_11_2  (
            .in0(_gnd_net_),
            .in1(N__36595),
            .in2(_gnd_net_),
            .in3(N__35184),
            .lcout(\PWMInstance2.periodCounterZ0Z_2 ),
            .ltout(),
            .carryin(\PWMInstance2.un1_periodCounter_2_cry_1 ),
            .carryout(\PWMInstance2.un1_periodCounter_2_cry_2 ),
            .clk(N__38677),
            .ce(),
            .sr(N__35310));
    defparam \PWMInstance2.periodCounter_3_LC_18_11_3 .C_ON=1'b1;
    defparam \PWMInstance2.periodCounter_3_LC_18_11_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.periodCounter_3_LC_18_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance2.periodCounter_3_LC_18_11_3  (
            .in0(_gnd_net_),
            .in1(N__35179),
            .in2(_gnd_net_),
            .in3(N__35163),
            .lcout(\PWMInstance2.periodCounterZ0Z_3 ),
            .ltout(),
            .carryin(\PWMInstance2.un1_periodCounter_2_cry_2 ),
            .carryout(\PWMInstance2.un1_periodCounter_2_cry_3 ),
            .clk(N__38677),
            .ce(),
            .sr(N__35310));
    defparam \PWMInstance2.periodCounter_4_LC_18_11_4 .C_ON=1'b1;
    defparam \PWMInstance2.periodCounter_4_LC_18_11_4 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.periodCounter_4_LC_18_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance2.periodCounter_4_LC_18_11_4  (
            .in0(_gnd_net_),
            .in1(N__36574),
            .in2(_gnd_net_),
            .in3(N__35160),
            .lcout(\PWMInstance2.periodCounterZ0Z_4 ),
            .ltout(),
            .carryin(\PWMInstance2.un1_periodCounter_2_cry_3 ),
            .carryout(\PWMInstance2.un1_periodCounter_2_cry_4 ),
            .clk(N__38677),
            .ce(),
            .sr(N__35310));
    defparam \PWMInstance2.periodCounter_5_LC_18_11_5 .C_ON=1'b1;
    defparam \PWMInstance2.periodCounter_5_LC_18_11_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.periodCounter_5_LC_18_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance2.periodCounter_5_LC_18_11_5  (
            .in0(_gnd_net_),
            .in1(N__35233),
            .in2(_gnd_net_),
            .in3(N__35157),
            .lcout(\PWMInstance2.periodCounterZ0Z_5 ),
            .ltout(),
            .carryin(\PWMInstance2.un1_periodCounter_2_cry_4 ),
            .carryout(\PWMInstance2.un1_periodCounter_2_cry_5 ),
            .clk(N__38677),
            .ce(),
            .sr(N__35310));
    defparam \PWMInstance2.periodCounter_6_LC_18_11_6 .C_ON=1'b1;
    defparam \PWMInstance2.periodCounter_6_LC_18_11_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.periodCounter_6_LC_18_11_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance2.periodCounter_6_LC_18_11_6  (
            .in0(_gnd_net_),
            .in1(N__35152),
            .in2(_gnd_net_),
            .in3(N__35133),
            .lcout(\PWMInstance2.periodCounterZ0Z_6 ),
            .ltout(),
            .carryin(\PWMInstance2.un1_periodCounter_2_cry_5 ),
            .carryout(\PWMInstance2.un1_periodCounter_2_cry_6 ),
            .clk(N__38677),
            .ce(),
            .sr(N__35310));
    defparam \PWMInstance2.periodCounter_7_LC_18_11_7 .C_ON=1'b1;
    defparam \PWMInstance2.periodCounter_7_LC_18_11_7 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.periodCounter_7_LC_18_11_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance2.periodCounter_7_LC_18_11_7  (
            .in0(N__35371),
            .in1(N__35130),
            .in2(_gnd_net_),
            .in3(N__35112),
            .lcout(\PWMInstance2.periodCounterZ0Z_7 ),
            .ltout(),
            .carryin(\PWMInstance2.un1_periodCounter_2_cry_6 ),
            .carryout(\PWMInstance2.un1_periodCounter_2_cry_7 ),
            .clk(N__38677),
            .ce(),
            .sr(N__35310));
    defparam \PWMInstance2.periodCounter_8_LC_18_12_0 .C_ON=1'b1;
    defparam \PWMInstance2.periodCounter_8_LC_18_12_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.periodCounter_8_LC_18_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance2.periodCounter_8_LC_18_12_0  (
            .in0(_gnd_net_),
            .in1(N__35108),
            .in2(_gnd_net_),
            .in3(N__35091),
            .lcout(\PWMInstance2.periodCounterZ0Z_8 ),
            .ltout(),
            .carryin(bfn_18_12_0_),
            .carryout(\PWMInstance2.un1_periodCounter_2_cry_8 ),
            .clk(N__38669),
            .ce(),
            .sr(N__35309));
    defparam \PWMInstance2.periodCounter_9_LC_18_12_1 .C_ON=1'b1;
    defparam \PWMInstance2.periodCounter_9_LC_18_12_1 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.periodCounter_9_LC_18_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance2.periodCounter_9_LC_18_12_1  (
            .in0(_gnd_net_),
            .in1(N__35457),
            .in2(_gnd_net_),
            .in3(N__35439),
            .lcout(\PWMInstance2.periodCounterZ0Z_9 ),
            .ltout(),
            .carryin(\PWMInstance2.un1_periodCounter_2_cry_8 ),
            .carryout(\PWMInstance2.un1_periodCounter_2_cry_9 ),
            .clk(N__38669),
            .ce(),
            .sr(N__35309));
    defparam \PWMInstance2.periodCounter_10_LC_18_12_2 .C_ON=1'b1;
    defparam \PWMInstance2.periodCounter_10_LC_18_12_2 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.periodCounter_10_LC_18_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance2.periodCounter_10_LC_18_12_2  (
            .in0(_gnd_net_),
            .in1(N__36217),
            .in2(_gnd_net_),
            .in3(N__35436),
            .lcout(\PWMInstance2.periodCounterZ0Z_10 ),
            .ltout(),
            .carryin(\PWMInstance2.un1_periodCounter_2_cry_9 ),
            .carryout(\PWMInstance2.un1_periodCounter_2_cry_10 ),
            .clk(N__38669),
            .ce(),
            .sr(N__35309));
    defparam \PWMInstance2.periodCounter_11_LC_18_12_3 .C_ON=1'b1;
    defparam \PWMInstance2.periodCounter_11_LC_18_12_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.periodCounter_11_LC_18_12_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance2.periodCounter_11_LC_18_12_3  (
            .in0(N__35369),
            .in1(N__36196),
            .in2(_gnd_net_),
            .in3(N__35433),
            .lcout(\PWMInstance2.periodCounterZ0Z_11 ),
            .ltout(),
            .carryin(\PWMInstance2.un1_periodCounter_2_cry_10 ),
            .carryout(\PWMInstance2.un1_periodCounter_2_cry_11 ),
            .clk(N__38669),
            .ce(),
            .sr(N__35309));
    defparam \PWMInstance2.periodCounter_12_LC_18_12_4 .C_ON=1'b1;
    defparam \PWMInstance2.periodCounter_12_LC_18_12_4 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.periodCounter_12_LC_18_12_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance2.periodCounter_12_LC_18_12_4  (
            .in0(N__35368),
            .in1(N__36557),
            .in2(_gnd_net_),
            .in3(N__35430),
            .lcout(\PWMInstance2.periodCounterZ0Z_12 ),
            .ltout(),
            .carryin(\PWMInstance2.un1_periodCounter_2_cry_11 ),
            .carryout(\PWMInstance2.un1_periodCounter_2_cry_12 ),
            .clk(N__38669),
            .ce(),
            .sr(N__35309));
    defparam \PWMInstance2.periodCounter_13_LC_18_12_5 .C_ON=1'b1;
    defparam \PWMInstance2.periodCounter_13_LC_18_12_5 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.periodCounter_13_LC_18_12_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance2.periodCounter_13_LC_18_12_5  (
            .in0(N__35370),
            .in1(N__35426),
            .in2(_gnd_net_),
            .in3(N__35406),
            .lcout(\PWMInstance2.periodCounterZ0Z_13 ),
            .ltout(),
            .carryin(\PWMInstance2.un1_periodCounter_2_cry_12 ),
            .carryout(\PWMInstance2.un1_periodCounter_2_cry_13 ),
            .clk(N__38669),
            .ce(),
            .sr(N__35309));
    defparam \PWMInstance2.periodCounter_14_LC_18_12_6 .C_ON=1'b1;
    defparam \PWMInstance2.periodCounter_14_LC_18_12_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.periodCounter_14_LC_18_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance2.periodCounter_14_LC_18_12_6  (
            .in0(_gnd_net_),
            .in1(N__36617),
            .in2(_gnd_net_),
            .in3(N__35403),
            .lcout(\PWMInstance2.periodCounterZ0Z_14 ),
            .ltout(),
            .carryin(\PWMInstance2.un1_periodCounter_2_cry_13 ),
            .carryout(\PWMInstance2.un1_periodCounter_2_cry_14 ),
            .clk(N__38669),
            .ce(),
            .sr(N__35309));
    defparam \PWMInstance2.periodCounter_15_LC_18_12_7 .C_ON=1'b1;
    defparam \PWMInstance2.periodCounter_15_LC_18_12_7 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.periodCounter_15_LC_18_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \PWMInstance2.periodCounter_15_LC_18_12_7  (
            .in0(_gnd_net_),
            .in1(N__35399),
            .in2(_gnd_net_),
            .in3(N__35379),
            .lcout(\PWMInstance2.periodCounterZ0Z_15 ),
            .ltout(),
            .carryin(\PWMInstance2.un1_periodCounter_2_cry_14 ),
            .carryout(\PWMInstance2.un1_periodCounter_2_cry_15 ),
            .clk(N__38669),
            .ce(),
            .sr(N__35309));
    defparam \PWMInstance2.periodCounter_16_LC_18_13_0 .C_ON=1'b0;
    defparam \PWMInstance2.periodCounter_16_LC_18_13_0 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.periodCounter_16_LC_18_13_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PWMInstance2.periodCounter_16_LC_18_13_0  (
            .in0(N__35372),
            .in1(N__35333),
            .in2(_gnd_net_),
            .in3(N__35337),
            .lcout(\PWMInstance2.periodCounterZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38657),
            .ce(),
            .sr(N__35308));
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_18_14_0 .C_ON=1'b0;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_18_14_0 .SEQ_MODE=4'b0000;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_18_14_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \PWMInstance2.un1_PWMPulseWidthCount_0_I_15_c_RNO_LC_18_14_0  (
            .in0(N__36575),
            .in1(N__36225),
            .in2(N__35238),
            .in3(N__36384),
            .lcout(\PWMInstance2.un1_PWMPulseWidthCount_0_I_15_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.periodCounter_RNIV91B_14_LC_18_14_1 .C_ON=1'b0;
    defparam \PWMInstance2.periodCounter_RNIV91B_14_LC_18_14_1 .SEQ_MODE=4'b0000;
    defparam \PWMInstance2.periodCounter_RNIV91B_14_LC_18_14_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \PWMInstance2.periodCounter_RNIV91B_14_LC_18_14_1  (
            .in0(_gnd_net_),
            .in1(N__36618),
            .in2(_gnd_net_),
            .in3(N__36596),
            .lcout(),
            .ltout(\PWMInstance2.un1_periodCounter12_1_0_a2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.periodCounter_RNI3BPO_10_LC_18_14_2 .C_ON=1'b0;
    defparam \PWMInstance2.periodCounter_RNI3BPO_10_LC_18_14_2 .SEQ_MODE=4'b0000;
    defparam \PWMInstance2.periodCounter_RNI3BPO_10_LC_18_14_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \PWMInstance2.periodCounter_RNI3BPO_10_LC_18_14_2  (
            .in0(N__36576),
            .in1(N__36558),
            .in2(N__36537),
            .in3(N__36219),
            .lcout(\PWMInstance2.un1_periodCounter12_1_0_a2_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.PWMPulseWidthCount_esr_4_LC_18_14_3 .C_ON=1'b0;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_4_LC_18_14_3 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_4_LC_18_14_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \PWMInstance2.PWMPulseWidthCount_esr_4_LC_18_14_3  (
            .in0(N__36501),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PWMInstance2.PWMPulseWidthCountZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38647),
            .ce(N__35865),
            .sr(N__35796));
    defparam \PWMInstance2.PWMPulseWidthCount_esr_5_LC_18_14_4 .C_ON=1'b0;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_5_LC_18_14_4 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_5_LC_18_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance2.PWMPulseWidthCount_esr_5_LC_18_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36345),
            .lcout(\PWMInstance2.PWMPulseWidthCountZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38647),
            .ce(N__35865),
            .sr(N__35796));
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_18_14_5 .C_ON=1'b0;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_18_14_5 .SEQ_MODE=4'b0000;
    defparam \PWMInstance2.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_18_14_5 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \PWMInstance2.un1_PWMPulseWidthCount_0_I_33_c_RNO_LC_18_14_5  (
            .in0(N__36218),
            .in1(N__35871),
            .in2(N__36201),
            .in3(N__36021),
            .lcout(\PWMInstance2.un1_PWMPulseWidthCount_0_I_33_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PWMInstance2.PWMPulseWidthCount_esr_10_LC_18_14_6 .C_ON=1'b0;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_10_LC_18_14_6 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_10_LC_18_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance2.PWMPulseWidthCount_esr_10_LC_18_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36150),
            .lcout(\PWMInstance2.PWMPulseWidthCountZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38647),
            .ce(N__35865),
            .sr(N__35796));
    defparam \PWMInstance2.PWMPulseWidthCount_esr_11_LC_18_14_7 .C_ON=1'b0;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_11_LC_18_14_7 .SEQ_MODE=4'b1000;
    defparam \PWMInstance2.PWMPulseWidthCount_esr_11_LC_18_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PWMInstance2.PWMPulseWidthCount_esr_11_LC_18_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36013),
            .lcout(\PWMInstance2.PWMPulseWidthCountZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38647),
            .ce(N__35865),
            .sr(N__35796));
    defparam PWM2_obufLegalizeSB_DFF_LC_18_20_0.C_ON=1'b0;
    defparam PWM2_obufLegalizeSB_DFF_LC_18_20_0.SEQ_MODE=4'b1000;
    defparam PWM2_obufLegalizeSB_DFF_LC_18_20_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 PWM2_obufLegalizeSB_DFF_LC_18_20_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PWM2_obufLegalizeSB_DFFNet),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36916),
            .ce(),
            .sr(_gnd_net_));
    defparam PWM3_obufLegalizeSB_DFF_LC_18_20_1.C_ON=1'b0;
    defparam PWM3_obufLegalizeSB_DFF_LC_18_20_1.SEQ_MODE=4'b1000;
    defparam PWM3_obufLegalizeSB_DFF_LC_18_20_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 PWM3_obufLegalizeSB_DFF_LC_18_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PWM3_obufLegalizeSB_DFFNet),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36916),
            .ce(),
            .sr(_gnd_net_));
    defparam MISO_obufLegalizeSB_DFF_LC_20_1_0.C_ON=1'b0;
    defparam MISO_obufLegalizeSB_DFF_LC_20_1_0.SEQ_MODE=4'b1000;
    defparam MISO_obufLegalizeSB_DFF_LC_20_1_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 MISO_obufLegalizeSB_DFF_LC_20_1_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(MISO_obufLegalizeSB_DFFNet),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__36906),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_2_5_LC_20_6_5.C_ON=1'b0;
    defparam OutReg_ess_RNO_2_5_LC_20_6_5.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_2_5_LC_20_6_5.LUT_INIT=16'b1100000010111011;
    LogicCell40 OutReg_ess_RNO_2_5_LC_20_6_5 (
            .in0(N__36873),
            .in1(N__38158),
            .in2(N__36831),
            .in3(N__36795),
            .lcout(OutReg_ess_RNO_2Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_1_5_LC_20_7_0.C_ON=1'b0;
    defparam OutReg_ess_RNO_1_5_LC_20_7_0.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_1_5_LC_20_7_0.LUT_INIT=16'b1000100011110011;
    LogicCell40 OutReg_ess_RNO_1_5_LC_20_7_0 (
            .in0(N__36783),
            .in1(N__37759),
            .in2(N__36750),
            .in3(N__36711),
            .lcout(),
            .ltout(OutReg_ess_RNO_1Z0Z_5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_0_5_LC_20_7_1.C_ON=1'b0;
    defparam OutReg_ess_RNO_0_5_LC_20_7_1.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_0_5_LC_20_7_1.LUT_INIT=16'b1111001111000000;
    LogicCell40 OutReg_ess_RNO_0_5_LC_20_7_1 (
            .in0(_gnd_net_),
            .in1(N__37565),
            .in2(N__36696),
            .in3(N__36693),
            .lcout(OutReg_ess_RNO_0Z0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_5_LC_20_8_0.C_ON=1'b0;
    defparam OutReg_ess_5_LC_20_8_0.SEQ_MODE=4'b1001;
    defparam OutReg_ess_5_LC_20_8_0.LUT_INIT=16'b1111000011100100;
    LogicCell40 OutReg_ess_5_LC_20_8_0 (
            .in0(N__38901),
            .in1(N__36687),
            .in2(N__36681),
            .in3(N__37387),
            .lcout(OutRegZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38714),
            .ce(N__37243),
            .sr(N__37137));
    defparam dataOut_RNO_0_LC_20_9_0.C_ON=1'b0;
    defparam dataOut_RNO_0_LC_20_9_0.SEQ_MODE=4'b0000;
    defparam dataOut_RNO_0_LC_20_9_0.LUT_INIT=16'b0101000001110011;
    LogicCell40 dataOut_RNO_0_LC_20_9_0 (
            .in0(N__39053),
            .in1(N__38864),
            .in2(N__39090),
            .in3(N__37344),
            .lcout(),
            .ltout(dataOut_RNOZ0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dataOut_LC_20_9_1.C_ON=1'b0;
    defparam dataOut_LC_20_9_1.SEQ_MODE=4'b1000;
    defparam dataOut_LC_20_9_1.LUT_INIT=16'b1100000011001010;
    LogicCell40 dataOut_LC_20_9_1 (
            .in0(N__36654),
            .in1(N__36629),
            .in2(N__36642),
            .in3(N__39056),
            .lcout(MISO_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38708),
            .ce(),
            .sr(_gnd_net_));
    defparam SSELr_0_LC_20_9_2.C_ON=1'b0;
    defparam SSELr_0_LC_20_9_2.SEQ_MODE=4'b1000;
    defparam SSELr_0_LC_20_9_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 SSELr_0_LC_20_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37863),
            .lcout(SSELrZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38708),
            .ce(),
            .sr(_gnd_net_));
    defparam bit_count_RNI8CK3_0_LC_20_9_3.C_ON=1'b0;
    defparam bit_count_RNI8CK3_0_LC_20_9_3.SEQ_MODE=4'b0000;
    defparam bit_count_RNI8CK3_0_LC_20_9_3.LUT_INIT=16'b0000000010001000;
    LogicCell40 bit_count_RNI8CK3_0_LC_20_9_3 (
            .in0(N__37810),
            .in1(N__38760),
            .in2(_gnd_net_),
            .in3(N__38798),
            .lcout(un1_bit_count_1_c1),
            .ltout(un1_bit_count_1_c1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam bit_count_2_LC_20_9_4.C_ON=1'b0;
    defparam bit_count_2_LC_20_9_4.SEQ_MODE=4'b1000;
    defparam bit_count_2_LC_20_9_4.LUT_INIT=16'b0001010101000000;
    LogicCell40 bit_count_2_LC_20_9_4 (
            .in0(N__39054),
            .in1(N__37887),
            .in2(N__37845),
            .in3(N__37962),
            .lcout(bit_countZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38708),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_ess_RNO_0_15_LC_20_9_5.C_ON=1'b0;
    defparam OutReg_ess_RNO_0_15_LC_20_9_5.SEQ_MODE=4'b0000;
    defparam OutReg_ess_RNO_0_15_LC_20_9_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 OutReg_ess_RNO_0_15_LC_20_9_5 (
            .in0(N__37564),
            .in1(N__37842),
            .in2(_gnd_net_),
            .in3(N__37830),
            .lcout(OutReg_ess_RNO_0Z0Z_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam bit_count_0_LC_20_9_7.C_ON=1'b0;
    defparam bit_count_0_LC_20_9_7.SEQ_MODE=4'b1000;
    defparam bit_count_0_LC_20_9_7.LUT_INIT=16'b0000000010100110;
    LogicCell40 bit_count_0_LC_20_9_7 (
            .in0(N__37811),
            .in1(N__38761),
            .in2(N__38805),
            .in3(N__39055),
            .lcout(bit_countZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38708),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_esr_RNO_1_8_LC_20_10_0.C_ON=1'b0;
    defparam OutReg_esr_RNO_1_8_LC_20_10_0.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_1_8_LC_20_10_0.LUT_INIT=16'b1000100011110011;
    LogicCell40 OutReg_esr_RNO_1_8_LC_20_10_0 (
            .in0(N__37794),
            .in1(N__37760),
            .in2(N__37617),
            .in3(N__37578),
            .lcout(),
            .ltout(OutReg_esr_RNO_1Z0Z_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_esr_RNO_0_8_LC_20_10_1.C_ON=1'b0;
    defparam OutReg_esr_RNO_0_8_LC_20_10_1.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_0_8_LC_20_10_1.LUT_INIT=16'b1111010110100000;
    LogicCell40 OutReg_esr_RNO_0_8_LC_20_10_1 (
            .in0(N__37569),
            .in1(_gnd_net_),
            .in2(N__37410),
            .in3(N__38001),
            .lcout(),
            .ltout(OutReg_esr_RNO_0Z0Z_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam OutReg_esr_8_LC_20_10_2.C_ON=1'b0;
    defparam OutReg_esr_8_LC_20_10_2.SEQ_MODE=4'b1000;
    defparam OutReg_esr_8_LC_20_10_2.LUT_INIT=16'b1010101010111000;
    LogicCell40 OutReg_esr_8_LC_20_10_2 (
            .in0(N__37407),
            .in1(N__38865),
            .in2(N__37398),
            .in3(N__37381),
            .lcout(OutRegZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38701),
            .ce(N__37240),
            .sr(N__37134));
    defparam OutReg_esr_RNO_2_8_LC_20_10_4.C_ON=1'b0;
    defparam OutReg_esr_RNO_2_8_LC_20_10_4.SEQ_MODE=4'b0000;
    defparam OutReg_esr_RNO_2_8_LC_20_10_4.LUT_INIT=16'b1010000011001111;
    LogicCell40 OutReg_esr_RNO_2_8_LC_20_10_4 (
            .in0(N__37017),
            .in1(N__36980),
            .in2(N__38166),
            .in3(N__38013),
            .lcout(OutReg_esr_RNO_2Z0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SSELr_1_LC_20_11_7.C_ON=1'b0;
    defparam SSELr_1_LC_20_11_7.SEQ_MODE=4'b1000;
    defparam SSELr_1_LC_20_11_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 SSELr_1_LC_20_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37995),
            .lcout(SSELrZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38694),
            .ce(),
            .sr(_gnd_net_));
    defparam SSELr_2_LC_20_12_6.C_ON=1'b0;
    defparam SSELr_2_LC_20_12_6.SEQ_MODE=4'b1000;
    defparam SSELr_2_LC_20_12_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 SSELr_2_LC_20_12_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39046),
            .lcout(SSELrZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38687),
            .ce(),
            .sr(_gnd_net_));
    defparam SCKr_0_LC_21_4_0.C_ON=1'b0;
    defparam SCKr_0_LC_21_4_0.SEQ_MODE=4'b1000;
    defparam SCKr_0_LC_21_4_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 SCKr_0_LC_21_4_0 (
            .in0(N__37971),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(SCKrZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38724),
            .ce(),
            .sr(_gnd_net_));
    defparam bit_count_RNI9MD6_2_LC_21_9_2.C_ON=1'b0;
    defparam bit_count_RNI9MD6_2_LC_21_9_2.SEQ_MODE=4'b0000;
    defparam bit_count_RNI9MD6_2_LC_21_9_2.LUT_INIT=16'b1000100000000000;
    LogicCell40 bit_count_RNI9MD6_2_LC_21_9_2 (
            .in0(N__37895),
            .in1(N__37960),
            .in2(_gnd_net_),
            .in3(N__37884),
            .lcout(un1_bit_count_1_c3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SCKr_RNIBA7C_2_LC_21_9_3.C_ON=1'b0;
    defparam SCKr_RNIBA7C_2_LC_21_9_3.SEQ_MODE=4'b0000;
    defparam SCKr_RNIBA7C_2_LC_21_9_3.LUT_INIT=16'b1000100010101010;
    LogicCell40 SCKr_RNIBA7C_2_LC_21_9_3 (
            .in0(N__39047),
            .in1(N__38758),
            .in2(_gnd_net_),
            .in3(N__38796),
            .lcout(SCKr_RNIBA7CZ0Z_2),
            .ltout(SCKr_RNIBA7CZ0Z_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SCKr_RNIMKEO_2_LC_21_9_4.C_ON=1'b0;
    defparam SCKr_RNIMKEO_2_LC_21_9_4.SEQ_MODE=4'b0000;
    defparam SCKr_RNIMKEO_2_LC_21_9_4.LUT_INIT=16'b1111111111110010;
    LogicCell40 SCKr_RNIMKEO_2_LC_21_9_4 (
            .in0(N__38797),
            .in1(N__38759),
            .in2(N__37926),
            .in3(N__39048),
            .lcout(N_45_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SCKr_1_LC_21_9_5.C_ON=1'b0;
    defparam SCKr_1_LC_21_9_5.SEQ_MODE=4'b1000;
    defparam SCKr_1_LC_21_9_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 SCKr_1_LC_21_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37905),
            .lcout(SCKrZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38715),
            .ce(),
            .sr(_gnd_net_));
    defparam bit_count_1_LC_21_9_6.C_ON=1'b0;
    defparam bit_count_1_LC_21_9_6.SEQ_MODE=4'b1000;
    defparam bit_count_1_LC_21_9_6.LUT_INIT=16'b0001000100100010;
    LogicCell40 bit_count_1_LC_21_9_6 (
            .in0(N__37896),
            .in1(N__39049),
            .in2(_gnd_net_),
            .in3(N__37885),
            .lcout(bit_countZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38715),
            .ce(),
            .sr(_gnd_net_));
    defparam bit_count_4_LC_21_10_2.C_ON=1'b0;
    defparam bit_count_4_LC_21_10_2.SEQ_MODE=4'b1000;
    defparam bit_count_4_LC_21_10_2.LUT_INIT=16'b0001001000100010;
    LogicCell40 bit_count_4_LC_21_10_2 (
            .in0(N__38967),
            .in1(N__39036),
            .in2(N__38997),
            .in3(N__38985),
            .lcout(bit_countZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38709),
            .ce(),
            .sr(_gnd_net_));
    defparam bit_count_RNIU615_0_4_LC_21_10_3.C_ON=1'b0;
    defparam bit_count_RNIU615_0_4_LC_21_10_3.SEQ_MODE=4'b0000;
    defparam bit_count_RNIU615_0_4_LC_21_10_3.LUT_INIT=16'b1100111111011111;
    LogicCell40 bit_count_RNIU615_0_4_LC_21_10_3 (
            .in0(N__38966),
            .in1(N__38794),
            .in2(N__38763),
            .in3(N__38983),
            .lcout(bit_count_RNIU615_0Z0Z_4),
            .ltout(bit_count_RNIU615_0Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SSELr_RNIGO0F_1_LC_21_10_4.C_ON=1'b0;
    defparam SSELr_RNIGO0F_1_LC_21_10_4.SEQ_MODE=4'b0000;
    defparam SSELr_RNIGO0F_1_LC_21_10_4.LUT_INIT=16'b0000000000001111;
    LogicCell40 SSELr_RNIGO0F_1_LC_21_10_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__39081),
            .in3(N__39034),
            .lcout(SSELr_RNIGO0FZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam bit_count_3_LC_21_10_5.C_ON=1'b0;
    defparam bit_count_3_LC_21_10_5.SEQ_MODE=4'b1000;
    defparam bit_count_3_LC_21_10_5.LUT_INIT=16'b0001000101000100;
    LogicCell40 bit_count_3_LC_21_10_5 (
            .in0(N__39035),
            .in1(N__38993),
            .in2(_gnd_net_),
            .in3(N__38984),
            .lcout(bit_countZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38709),
            .ce(),
            .sr(_gnd_net_));
    defparam bit_count_RNIU615_4_LC_21_10_6.C_ON=1'b0;
    defparam bit_count_RNIU615_4_LC_21_10_6.SEQ_MODE=4'b0000;
    defparam bit_count_RNIU615_4_LC_21_10_6.LUT_INIT=16'b1111111011111111;
    LogicCell40 bit_count_RNIU615_4_LC_21_10_6 (
            .in0(N__38982),
            .in1(N__38965),
            .in2(N__38762),
            .in3(N__38793),
            .lcout(un1_OutReg51_4_0_i_o3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SCKr_2_LC_21_10_7.C_ON=1'b0;
    defparam SCKr_2_LC_21_10_7.SEQ_MODE=4'b1000;
    defparam SCKr_2_LC_21_10_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 SCKr_2_LC_21_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38795),
            .lcout(SCKrZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38709),
            .ce(),
            .sr(_gnd_net_));
endmodule // SPI
